----------------------------------------------------------------------------------
--                            Tabla de nombre                                   --
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library WORK;
use WORK.VGA_PKG.ALL;

entity tabla_nombre is
	port (
	--Puertos de entrada
	clk          	  : in std_logic;
	dir_tabla_nombre  : in std_logic_vector(10-1 downto 0); --960 posiciones de memoria
 	--Puertos de salida
	dato_tabla_nombre : out std_logic_vector(8-1 downto 0)
);
end tabla_nombre;

architecture behavioral of tabla_nombre is

signal dir_int_img : natural range 0 to 2**10-1;
type img is array (natural range<>) of std_logic_vector(8-1 downto 0);
constant title : img := (
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00010110",
	"00001010",
	"00011011",
	"00010010",
	"00011000",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100000",
	"00011000",
	"00011011",
	"00010101",
	"00001101",
	"00100100",
	"00100100",
	"00011101",
	"00010010",
	"00010110",
	"00001110",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00110110",
	"00110111",
	"00110110",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00110101",
	"00100101",
	"00100101",
	"00100101",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00110110",
	"00110111",
	"00110110",
	"00110111",
	"00110110",
	"00110111",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00111001",
	"00111010",
	"00111011",
	"00111010",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00110101",
	"00100101",
	"00100101",
	"00100101",
	"00100101",
	"00100101",
	"00100101",
	"00111000",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00111001",
	"00111010",
	"00111011",
	"00111010",
	"00111011",
	"00111010",
	"00111011",
	"00111100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"01000101",
	"01000101",
	"01000101",
	"01000101",
	"01000101",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"01000101",
	"01000101",
	"01010011",
	"01010100",
	"01010011",
	"01010100",
	"01000101",
	"01000101",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"01000111",
	"01000111",
	"01000111",
	"01000111",
	"01000111",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"01000111",
	"01000111",
	"01010101",
	"01010110",
	"01010101",
	"01010110",
	"01000111",
	"01000111",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"01000101",
	"01000101",
	"01000101",
	"01000101",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"01000111",
	"01000111",
	"01000111",
	"01000111",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00110110",
	"00110111",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00110101",
	"00100101",
	"00100101",
	"00111000",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"00100100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110101",
	"10110100",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110",
	"10110111",
	"10110110"
);

begin

dir_int_img <= to_integer(unsigned(dir_tabla_nombre));

P_img: process (clk)
begin
	if clk'event and clk='1' then
		dato_tabla_nombre <= title(dir_int_img);
	end if;
end process;

end behavioral;