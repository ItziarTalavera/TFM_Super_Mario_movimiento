----------------------------------------------------------------------------------
--                              Tabla patrones                                  --
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library WORK;
use WORK.VGA_PKG.ALL;

entity tabla_patrones is
port(
	--Puertos de entrada
	clk                 : in std_logic;
	dir_tabla_patrones  : in std_logic_vector(13-1 downto 0); --8192 posiciones de memoria (8 KiB)
 	--Puertos de salida
	dato_tabla_patrones : out std_logic_vector(8-1 downto 0)
);
end tabla_patrones;

architecture behavioral of tabla_patrones is

signal dir_int_img : natural range 0 to 2**13-1;
type img is array (natural range<>) of std_logic_vector (8-1 downto 0);
constant title : img := (
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00011100",
	"00110010",
	"01100011",
	"01100011",
	"01100011",
	"00100110",
	"00011100",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00011000",
	"00011100",
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"01111110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00111110",
	"01100011",
	"01110000",
	"00111100",
	"00011110",
	"00000111",
	"01111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01111110",
	"00110000",
	"00011000",
	"00111100",
	"01100000",
	"01100011",
	"00111110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00111000",
	"00111100",
	"00110110",
	"00110011",
	"01111111",
	"00110000",
	"00110000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00111111",
	"00000011",
	"00111111",
	"01100000",
	"01100000",
	"01100011",
	"00111110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00111100",
	"00000110",
	"00000011",
	"00111111",
	"01100011",
	"01100011",
	"00111110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01111111",
	"01100011",
	"00110000",
	"00011000",
	"00001100",
	"00001100",
	"00001100",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00111110",
	"01100011",
	"01100011",
	"00111110",
	"01100011",
	"01100011",
	"00111110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00111110",
	"01100011",
	"01100011",
	"01111110",
	"01100000",
	"00110000",
	"00011110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00011100",
	"00110110",
	"01100011",
	"01100011",
	"01111111",
	"01100011",
	"01100011",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00111111",
	"01100011",
	"01100011",
	"00111111",
	"01100011",
	"01100011",
	"00111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00111100",
	"01100110",
	"00000011",
	"00000011",
	"00000011",
	"01100110",
	"00111100",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00011111",
	"00110011",
	"01100011",
	"01100011",
	"01100011",
	"00110011",
	"00011111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01111111",
	"00000011",
	"00000011",
	"00111111",
	"00000011",
	"00000011",
	"01111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01111111",
	"00000011",
	"00000011",
	"00111111",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01111100",
	"00000110",
	"00000011",
	"01110011",
	"01100011",
	"01100110",
	"01111100",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01100011",
	"01100011",
	"01100011",
	"01111111",
	"01100011",
	"01100011",
	"01100011",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01111110",
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"01111110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01111000",
	"01100000",
	"01100000",
	"01100000",
	"01100011",
	"01100011",
	"00111110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01100011",
	"00110011",
	"00011011",
	"00001111",
	"00011111",
	"00111011",
	"01110011",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000110",
	"00000110",
	"00000110",
	"00000110",
	"00000110",
	"00000110",
	"01111110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01100011",
	"01110111",
	"01111111",
	"01111111",
	"01101011",
	"01100011",
	"01100011",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01100011",
	"01100111",
	"01101111",
	"01111111",
	"01111011",
	"01110011",
	"01100011",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00111110",
	"01100011",
	"01100011",
	"01100011",
	"01100011",
	"01100011",
	"00111110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00111111",
	"01100011",
	"01100011",
	"01100011",
	"00111111",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00111110",
	"01100011",
	"01100011",
	"01100011",
	"01111011",
	"00110011",
	"01011110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00111111",
	"01100011",
	"01100011",
	"01110011",
	"00011111",
	"00111011",
	"01110011",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00011110",
	"00110011",
	"00000011",
	"00111110",
	"01100000",
	"01100011",
	"00111110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01111110",
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01100011",
	"01100011",
	"01100011",
	"01100011",
	"01100011",
	"01100011",
	"00111110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01100011",
	"01100011",
	"01100011",
	"01110111",
	"00111110",
	"00011100",
	"00001000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01100011",
	"01100011",
	"01101011",
	"01111111",
	"01111111",
	"01110111",
	"01100011",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01100011",
	"01110111",
	"00111110",
	"00011100",
	"00111110",
	"01110111",
	"01100011",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01100110",
	"01100110",
	"01100110",
	"00111100",
	"00011000",
	"00011000",
	"00011000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01111111",
	"01110000",
	"00111000",
	"00011100",
	"00001110",
	"00000111",
	"01111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01111110",
	"01111110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00100010",
	"00010100",
	"00001000",
	"00010100",
	"00100010",
	"00000000",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00011000",
	"00111100",
	"00111100",
	"00111100",
	"00011000",
	"00011000",
	"00000000",
	"00011000",
	"11111111",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000000",
	"00111000",
	"01111100",
	"11111111",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111111",
	"11000111",
	"10000011",
	"11111110",
	"11111110",
	"11111110",
	"01111100",
	"00111000",
	"00000000",
	"00000000",
	"11111111",
	"00000001",
	"00000001",
	"00000001",
	"10000011",
	"11000111",
	"11111111",
	"11111111",
	"11111111",
	"00010000",
	"00100000",
	"00100000",
	"00100000",
	"00100000",
	"00100000",
	"00010000",
	"00000000",
	"00011100",
	"00111110",
	"00111110",
	"00111110",
	"00111110",
	"00111110",
	"00011100",
	"00000000",
	"11000000",
	"10100000",
	"11010000",
	"11010000",
	"11110000",
	"11110000",
	"11100000",
	"11000000",
	"11000000",
	"01100000",
	"00110000",
	"00110000",
	"00010000",
	"00010000",
	"00100000",
	"11000000",
	"10000000",
	"11000000",
	"11100000",
	"11110000",
	"11111000",
	"11111100",
	"11111110",
	"11111111",
	"10000000",
	"01000000",
	"00100000",
	"00010000",
	"00001000",
	"00000100",
	"00000010",
	"00000001",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11100000",
	"11111100",
	"11111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11100000",
	"00011100",
	"00000011",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000111",
	"00111111",
	"11111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000111",
	"00111000",
	"11000000",
	"00000001",
	"00000011",
	"00000111",
	"00001111",
	"00011111",
	"00111111",
	"01111111",
	"11111111",
	"00000001",
	"00000010",
	"00000100",
	"00001000",
	"00010000",
	"00100000",
	"01000000",
	"10000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00100000",
	"01110000",
	"01110000",
	"01110000",
	"01110110",
	"00100110",
	"00000110",
	"00000110",
	"11100000",
	"00010000",
	"00001000",
	"00000000",
	"00000110",
	"00000001",
	"00000001",
	"00000010",
	"11100000",
	"11110000",
	"11111000",
	"11111000",
	"11111110",
	"11111111",
	"11111111",
	"11111110",
	"11000000",
	"00100000",
	"00011000",
	"00000100",
	"00000100",
	"00000100",
	"01100010",
	"00010001",
	"11000000",
	"11100000",
	"11111000",
	"11111100",
	"11111100",
	"11111100",
	"10011110",
	"11101111",
	"00000011",
	"00000100",
	"00001000",
	"00101000",
	"01010000",
	"10000010",
	"10000100",
	"10000000",
	"00000011",
	"00000111",
	"00001111",
	"00101111",
	"01111111",
	"11111101",
	"11111011",
	"11111111",
	"00001001",
	"00010101",
	"00010010",
	"01010000",
	"10100000",
	"10000000",
	"10000000",
	"01000000",
	"00001001",
	"00011101",
	"00011111",
	"01011111",
	"11111111",
	"11111111",
	"11111111",
	"01111111",
	"00100100",
	"01001000",
	"10010000",
	"00010000",
	"11100000",
	"00000000",
	"00000000",
	"00000000",
	"11011100",
	"10111000",
	"01110000",
	"11110000",
	"11100000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000010",
	"11000111",
	"11111100",
	"00110000",
	"10000001",
	"01000110",
	"00111000",
	"11111111",
	"11111101",
	"00111000",
	"00000011",
	"11001111",
	"11111111",
	"01111110",
	"00111000",
	"00000010",
	"00000001",
	"01000011",
	"00111110",
	"00011100",
	"00000000",
	"11000011",
	"00111100",
	"11111101",
	"11111110",
	"10111100",
	"11000001",
	"11100011",
	"11111111",
	"11111111",
	"00111100",
	"00100000",
	"01000000",
	"10000000",
	"00000000",
	"01100000",
	"00011001",
	"00000110",
	"00000000",
	"00111111",
	"01111111",
	"11111111",
	"01111111",
	"01111111",
	"00011111",
	"00000110",
	"00000000",
	"00000011",
	"00000111",
	"00001111",
	"00001111",
	"00001111",
	"00001111",
	"00000111",
	"00000011",
	"00000011",
	"00000100",
	"00001000",
	"00001000",
	"00001000",
	"00001000",
	"00000100",
	"00000011",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00111000",
	"01111100",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111100",
	"11111110",
	"00000111",
	"00000011",
	"11111110",
	"11111110",
	"11111110",
	"01111100",
	"00111000",
	"00000000",
	"00000000",
	"00000000",
	"00010001",
	"00111001",
	"00010001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"01111111",
	"01111111",
	"01111111",
	"01111111",
	"01111111",
	"01111111",
	"01111111",
	"01111111",
	"00000000",
	"00010000",
	"00011000",
	"00011100",
	"00111111",
	"11111101",
	"01111010",
	"10011011",
	"00010000",
	"00101000",
	"00100100",
	"00100011",
	"11000000",
	"00000010",
	"10000101",
	"01100100",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00000000",
	"11111110",
	"11111110",
	"11100110",
	"11100110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"00000001",
	"00000001",
	"00011001",
	"00111001",
	"00110001",
	"00000001",
	"00000001",
	"00000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"10000000",
	"10000000",
	"11111111",
	"00001000",
	"00001000",
	"00001000",
	"11111111",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"10000000",
	"10000000",
	"10000000",
	"11111111",
	"00001000",
	"00001000",
	"00001000",
	"11111111",
	"00000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111111",
	"11111111",
	"11100111",
	"11100111",
	"11111111",
	"11111111",
	"11111111",
	"01111111",
	"10000000",
	"10000000",
	"10011000",
	"10111000",
	"10110000",
	"10000000",
	"10000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"11111100",
	"00000110",
	"00000010",
	"00000011",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"11111100",
	"11111110",
	"11111110",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"10000001",
	"01000010",
	"00111100",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"01111110",
	"00111100",
	"11111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"10000000",
	"01000001",
	"00111110",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"01111111",
	"00111110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"10000000",
	"11000001",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"01111111",
	"00111110",
	"00011111",
	"00100000",
	"01000000",
	"01000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"00011111",
	"00111111",
	"01111111",
	"01111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000001",
	"01000010",
	"00111100",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"01111110",
	"00111100",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00000000",
	"00010000",
	"00010000",
	"00010000",
	"00001000",
	"00001000",
	"00001000",
	"00000000",
	"11111110",
	"00000001",
	"00000101",
	"11100001",
	"11110001",
	"01110001",
	"01110001",
	"01100001",
	"00000000",
	"11111110",
	"11111110",
	"00011110",
	"11001110",
	"11001110",
	"11001110",
	"11111110",
	"01111111",
	"10000000",
	"10100000",
	"10000011",
	"10000111",
	"10001110",
	"10001110",
	"10001111",
	"00000000",
	"11111111",
	"11111111",
	"11111100",
	"11111001",
	"11111001",
	"11111001",
	"11111000",
	"10000001",
	"10000001",
	"00000001",
	"10000001",
	"10000001",
	"00000101",
	"00000001",
	"11111111",
	"01111110",
	"01111110",
	"11111110",
	"01111110",
	"01111110",
	"11111110",
	"11111110",
	"11111111",
	"10001111",
	"10000011",
	"10000011",
	"10000001",
	"10000011",
	"10100011",
	"10000000",
	"11111111",
	"11111110",
	"11111110",
	"11111111",
	"11111110",
	"11111110",
	"11111111",
	"11111111",
	"11111111",
	"11111110",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111110",
	"00000001",
	"00000101",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"01111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"01111111",
	"10000000",
	"10100000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111110",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000101",
	"00000001",
	"11111110",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"01111111",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10100000",
	"10000000",
	"01111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00011100",
	"00111110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00111111",
	"01111111",
	"11100000",
	"11000000",
	"01111111",
	"01111111",
	"01111111",
	"00111110",
	"00011100",
	"00000000",
	"00000000",
	"00000000",
	"10001000",
	"10011100",
	"10001000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"00000100",
	"11100111",
	"11100111",
	"11100111",
	"11100111",
	"11100111",
	"11110111",
	"00000000",
	"11110111",
	"00010100",
	"00010100",
	"00010100",
	"00010100",
	"00010100",
	"11110111",
	"00000000",
	"01000000",
	"01111110",
	"01111110",
	"01111110",
	"01111110",
	"01111110",
	"01111111",
	"00000000",
	"01111111",
	"01000001",
	"01000001",
	"01000001",
	"01000001",
	"01000001",
	"01111111",
	"00000000",
	"11111110",
	"11111110",
	"11111110",
	"11100110",
	"11100110",
	"11111110",
	"11111110",
	"11111110",
	"00000001",
	"00000001",
	"00000001",
	"00011001",
	"00111001",
	"00110001",
	"00000001",
	"11111110",
	"11111111",
	"00000001",
	"00111111",
	"00110001",
	"00110001",
	"00110001",
	"00110001",
	"00110001",
	"11111111",
	"11111111",
	"11000001",
	"11001111",
	"11001111",
	"11001111",
	"11001111",
	"11001111",
	"11111111",
	"00000000",
	"11110000",
	"10010000",
	"10010000",
	"10010000",
	"10010000",
	"10010000",
	"11111111",
	"11111111",
	"00001111",
	"01101111",
	"01101111",
	"01101111",
	"01101111",
	"01101111",
	"11111111",
	"00000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111111",
	"10000000",
	"11111111",
	"10010101",
	"10001011",
	"10010101",
	"10001011",
	"10010101",
	"11111111",
	"11111111",
	"10000000",
	"11101010",
	"11110100",
	"11101010",
	"11110100",
	"11101010",
	"00110001",
	"00110001",
	"00110001",
	"00110001",
	"00110001",
	"00110001",
	"11111111",
	"11111100",
	"11001111",
	"11001111",
	"11001111",
	"11001111",
	"11001111",
	"11001111",
	"11111111",
	"11111100",
	"10010000",
	"10010000",
	"10010000",
	"10010000",
	"10010000",
	"10010000",
	"11111111",
	"11111111",
	"01101111",
	"01101111",
	"01101111",
	"01101111",
	"01101111",
	"01101111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111111",
	"11111111",
	"10001011",
	"10010101",
	"10001011",
	"10010101",
	"10001011",
	"10010101",
	"11111111",
	"00111111",
	"11110100",
	"11101010",
	"11110100",
	"11101010",
	"11110100",
	"11101010",
	"11111111",
	"00111111",
	"11000100",
	"11000100",
	"11000100",
	"11000100",
	"11000100",
	"11000100",
	"11000100",
	"11000100",
	"00111100",
	"00111100",
	"00111100",
	"00111100",
	"00111100",
	"00111100",
	"00111100",
	"00111100",
	"00100000",
	"00100000",
	"00100000",
	"00100000",
	"00100000",
	"00100000",
	"00100000",
	"00100000",
	"11011111",
	"11011111",
	"11011111",
	"11011111",
	"11011111",
	"11011111",
	"11011111",
	"11011111",
	"00100010",
	"00100101",
	"00100010",
	"00100101",
	"00100010",
	"00100101",
	"00100010",
	"00100101",
	"00111101",
	"00111010",
	"00111101",
	"00111010",
	"00111101",
	"00111010",
	"00111101",
	"00111010",
	"11111000",
	"11111100",
	"11111110",
	"11111110",
	"11111111",
	"11111111",
	"11111111",
	"01111111",
	"11111000",
	"00000100",
	"00000010",
	"00000010",
	"00000001",
	"00000001",
	"00000001",
	"10000001",
	"11111111",
	"11111110",
	"11111110",
	"11111100",
	"00000000",
	"00000000",
	"10000000",
	"10000000",
	"11111111",
	"00000001",
	"00000001",
	"00000011",
	"11111111",
	"11111111",
	"01111111",
	"01111111",
	"11111111",
	"00000001",
	"00000001",
	"00000000",
	"00000000",
	"00011111",
	"00111111",
	"00111111",
	"11111111",
	"11111110",
	"11111110",
	"11111111",
	"11111111",
	"11100000",
	"11000000",
	"11000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"01111110",
	"00111100",
	"00000000",
	"11111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"10000001",
	"11000011",
	"11111111",
	"00011111",
	"00100000",
	"01000000",
	"01000000",
	"10111000",
	"11111100",
	"11111110",
	"11111110",
	"00011111",
	"00111111",
	"01111111",
	"01111111",
	"11000111",
	"10000011",
	"10000001",
	"10000001",
	"00111111",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000110",
	"11111000",
	"11000001",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111110",
	"11111000",
	"11000000",
	"11000000",
	"11000000",
	"11000000",
	"10000000",
	"10000000",
	"00000000",
	"11111111",
	"00111111",
	"00111111",
	"00111111",
	"00111111",
	"01111111",
	"01111111",
	"11111111",
	"11111111",
	"01111111",
	"01111111",
	"01111111",
	"01111111",
	"00111111",
	"00111111",
	"00011111",
	"11111111",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"11000000",
	"11000000",
	"11100000",
	"11111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111110",
	"11111100",
	"10111000",
	"10000000",
	"10000000",
	"10000000",
	"11000000",
	"01111111",
	"10000001",
	"10000011",
	"11000111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"01111111",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00100001",
	"01010011",
	"10001101",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11011111",
	"10101101",
	"01110011",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000100",
	"11001010",
	"10110001",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111011",
	"10110101",
	"11001110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11101110",
	"11111111",
	"11111111",
	"11111111",
	"11101110",
	"11101110",
	"11101110",
	"11101110",
	"11101110",
	"11101110",
	"11101110",
	"11101110",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11101110",
	"11101110",
	"11101110",
	"11101110",
	"11101110",
	"11101110",
	"11101110",
	"11101110",
	"11101110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111111",
	"11111111",
	"11111111",
	"11100111",
	"11100111",
	"11111111",
	"11111111",
	"01111111",
	"10000000",
	"10000000",
	"10000000",
	"10011000",
	"10111000",
	"10110000",
	"10000000",
	"01111111",
	"00000000",
	"10000100",
	"10000100",
	"10000010",
	"10000010",
	"10000010",
	"10000010",
	"10000010",
	"00000100",
	"00011110",
	"11111110",
	"01111111",
	"01111111",
	"01111111",
	"01111111",
	"01111111",
	"00000000",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00100000",
	"01011001",
	"01011111",
	"10111111",
	"10111111",
	"10111111",
	"10111111",
	"10111111",
	"10000100",
	"10000100",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"01111110",
	"00011100",
	"10000100",
	"00000000",
	"10000000",
	"00000000",
	"10000000",
	"00000000",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"01011111",
	"01010001",
	"00100001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"10000000",
	"10000000",
	"01100000",
	"00010000",
	"00011000",
	"00000100",
	"00000100",
	"00000011",
	"01000000",
	"00100000",
	"00000000",
	"00001000",
	"00000000",
	"00000010",
	"00000001",
	"00000000",
	"00100000",
	"00100000",
	"00100011",
	"00101111",
	"00101111",
	"00100000",
	"00100000",
	"10100000",
	"11010000",
	"11010000",
	"11011100",
	"11010000",
	"11011111",
	"11010000",
	"11010000",
	"01010000",
	"00001110",
	"00001111",
	"00001111",
	"11111111",
	"11111111",
	"00001111",
	"00001111",
	"00001110",
	"00001001",
	"00001000",
	"11111000",
	"00001000",
	"11111000",
	"00001000",
	"00001000",
	"00001001",
	"00000011",
	"11100001",
	"00011000",
	"00001101",
	"11100111",
	"11100111",
	"11110111",
	"11110111",
	"11111100",
	"00011110",
	"11100111",
	"11110011",
	"00011010",
	"00011010",
	"00001010",
	"00001001",
	"11110110",
	"11000010",
	"10111010",
	"11111100",
	"11111100",
	"11111110",
	"11111110",
	"11111111",
	"00001101",
	"00111111",
	"01000111",
	"10000011",
	"10000011",
	"11000001",
	"11110001",
	"01111110",
	"11000000",
	"11111111",
	"10001111",
	"01110110",
	"11110011",
	"11111011",
	"11111111",
	"11111111",
	"01111111",
	"11000000",
	"11110000",
	"10001001",
	"00001110",
	"00000110",
	"00000100",
	"10001100",
	"10111111",
	"11011111",
	"11011111",
	"11101111",
	"11101111",
	"11110000",
	"11111110",
	"11111111",
	"11111100",
	"11111100",
	"10111000",
	"10011100",
	"11011110",
	"11001111",
	"01100001",
	"01111111",
	"11111111",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"11111111",
	"11111111",
	"00000001",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00000001",
	"00000001",
	"11111111",
	"01111111",
	"11000000",
	"11000000",
	"11000000",
	"11000000",
	"11111111",
	"11111111",
	"11000000",
	"01111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11000000",
	"11000000",
	"11111111",
	"00000000",
	"11111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111111",
	"11111111",
	"00000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00000000",
	"00000000",
	"11000100",
	"11001111",
	"11010000",
	"11010000",
	"11010000",
	"11100000",
	"11111111",
	"11111111",
	"00111100",
	"00111111",
	"00111111",
	"00111111",
	"00111111",
	"00111111",
	"00100000",
	"00100000",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"11111111",
	"00000001",
	"00000001",
	"00000001",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00000001",
	"11111111",
	"11111111",
	"11111111",
	"11000000",
	"11000000",
	"11000000",
	"11000000",
	"11111111",
	"11000000",
	"11000000",
	"11000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11000000",
	"11111111",
	"11111111",
	"11111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111111",
	"00000000",
	"00000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00000000",
	"11111111",
	"11111111",
	"11100000",
	"11100000",
	"11000000",
	"11000000",
	"11000000",
	"11111111",
	"11000000",
	"11000000",
	"00111111",
	"00111111",
	"01111111",
	"01111111",
	"01111111",
	"01000000",
	"01111111",
	"01111111",
	"00000001",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"11000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11000000",
	"11000000",
	"11000000",
	"11000000",
	"11000000",
	"11000000",
	"11000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"01000000",
	"01000000",
	"01000000",
	"01000000",
	"01000000",
	"01000000",
	"00100000",
	"00100000",
	"11111111",
	"11111111",
	"10101011",
	"01010101",
	"10101011",
	"00000001",
	"00000001",
	"11111111",
	"00000001",
	"00000001",
	"01010101",
	"10101011",
	"01010101",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11101010",
	"11010101",
	"11101010",
	"11000000",
	"11000000",
	"01111111",
	"11000000",
	"11000000",
	"11010101",
	"11101010",
	"11010101",
	"11111111",
	"11111111",
	"01111111",
	"11111111",
	"01010101",
	"10101010",
	"01010101",
	"00000000",
	"00000000",
	"11111111",
	"00000000",
	"00000000",
	"10101010",
	"01010101",
	"10101010",
	"11111111",
	"11111111",
	"11111111",
	"00000000",
	"11111111",
	"11110101",
	"11101010",
	"11010101",
	"11010000",
	"11010000",
	"11001111",
	"11000100",
	"00100000",
	"00101010",
	"00110101",
	"00111010",
	"00111111",
	"00111111",
	"00111111",
	"00111100",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111100",
	"11111100",
	"11111100",
	"11111100",
	"00000000",
	"00000000",
	"00000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"01111110",
	"00111110",
	"00111110",
	"00011110",
	"00000000",
	"00000000",
	"00000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111000",
	"11110000",
	"11110000",
	"11100000",
	"00000000",
	"00000000",
	"00000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"01111111",
	"00111111",
	"00111111",
	"00011111",
	"00000000",
	"00000000",
	"00000000",
	"11111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111111",
	"11111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11100000",
	"11111000",
	"11111100",
	"11111111",
	"11111110",
	"11111110",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"10000111",
	"10011111",
	"10111111",
	"11111111",
	"01111111",
	"01111111",
	"11111111",
	"11111111",
	"00000000",
	"00000111",
	"00000111",
	"00000111",
	"00000111",
	"00000111",
	"00000111",
	"00000111",
	"00001111",
	"00001000",
	"00001000",
	"00001000",
	"00001000",
	"00001000",
	"00001000",
	"11111111",
	"00000000",
	"11110000",
	"11110000",
	"11110000",
	"11110000",
	"11110000",
	"11110000",
	"11110000",
	"11111000",
	"00001000",
	"00001000",
	"00001000",
	"00001000",
	"00001000",
	"00001000",
	"11111111",
	"00010010",
	"00010010",
	"00110110",
	"00000000",
	"00000000",
	"00000000",
	"01111111",
	"00000000",
	"01001001",
	"01001001",
	"01001001",
	"01111111",
	"01111111",
	"00000000",
	"00000000",
	"00000000",
	"10100000",
	"10100000",
	"10100011",
	"10101111",
	"00101111",
	"00100000",
	"00100000",
	"00100000",
	"01010000",
	"01010000",
	"01011100",
	"01010000",
	"11011111",
	"11010000",
	"11010000",
	"11010000",
	"00001110",
	"00001110",
	"00001110",
	"11111110",
	"11111110",
	"00001110",
	"00001110",
	"00001110",
	"00001001",
	"00001001",
	"11111001",
	"00001001",
	"11111001",
	"00001001",
	"00001001",
	"00001001",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"01111111",
	"01111101",
	"01110011",
	"00010000",
	"00010001",
	"10001001",
	"10001011",
	"11001010",
	"11001010",
	"11001110",
	"11111100",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11000000",
	"00100000",
	"00100000",
	"00100000",
	"00000000",
	"00000000",
	"11100000",
	"11110000",
	"00110000",
	"11011000",
	"11011000",
	"11011000",
	"00000000",
	"00000000",
	"00000110",
	"00001100",
	"00001100",
	"00011001",
	"00011001",
	"00011001",
	"00000000",
	"00000000",
	"00000111",
	"00001111",
	"00001111",
	"00011111",
	"00011111",
	"00011111",
	"00100000",
	"00100000",
	"00100000",
	"00100000",
	"00100000",
	"11000000",
	"00000000",
	"00000000",
	"11011000",
	"11011000",
	"11011000",
	"11011000",
	"11011000",
	"11110000",
	"11110000",
	"11100000",
	"00011001",
	"00011001",
	"00011001",
	"00011001",
	"00011001",
	"00001100",
	"00001100",
	"00000110",
	"00011111",
	"00011111",
	"00011111",
	"00011111",
	"00011111",
	"00001111",
	"00001111",
	"00000111",
	"11110000",
	"11110111",
	"11110111",
	"11110111",
	"11110111",
	"11110111",
	"11110111",
	"00000111",
	"10001111",
	"10001000",
	"10001000",
	"11111000",
	"00001000",
	"00001000",
	"00001000",
	"11111111",
	"00000111",
	"11110111",
	"11110111",
	"11110111",
	"11110111",
	"11110111",
	"11110111",
	"11110000",
	"11111000",
	"00001000",
	"00001000",
	"00001111",
	"00001000",
	"00001000",
	"00001000",
	"11111111",
	"00000001",
	"00000010",
	"00000100",
	"00001000",
	"11110000",
	"11110000",
	"11110000",
	"11110000",
	"11111110",
	"11111101",
	"11111011",
	"11110111",
	"00001111",
	"00001111",
	"00001111",
	"00001111",
	"11110000",
	"11110000",
	"11110000",
	"11110000",
	"11111000",
	"11111100",
	"11111110",
	"11111111",
	"00001111",
	"00001111",
	"00001111",
	"00001111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"10000000",
	"11000000",
	"11100000",
	"11110000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11110000",
	"11110000",
	"11110000",
	"11110000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11110000",
	"11110000",
	"11110000",
	"11110000",
	"11101111",
	"11011111",
	"10111111",
	"01111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00011000",
	"00011000",
	"11111000",
	"00000100",
	"00000010",
	"00000010",
	"00000010",
	"00000001",
	"01000001",
	"01000001",
	"11111000",
	"11111100",
	"11111110",
	"11111110",
	"11111110",
	"11111111",
	"11111111",
	"11111111",
	"01000001",
	"00000001",
	"00000101",
	"00100010",
	"11000010",
	"00000010",
	"10000100",
	"01111000",
	"11111111",
	"11111111",
	"11111111",
	"11111110",
	"11111110",
	"11111110",
	"11111100",
	"01111000",
	"00011111",
	"00100000",
	"01000000",
	"01000000",
	"01000000",
	"10000000",
	"10000010",
	"10000010",
	"00011111",
	"00111111",
	"01111111",
	"01111111",
	"01111111",
	"11111111",
	"11111111",
	"11111111",
	"10000010",
	"10000000",
	"10100000",
	"01000100",
	"01000011",
	"01000000",
	"00100001",
	"00011110",
	"11111111",
	"11111111",
	"11111111",
	"01111111",
	"01111111",
	"01111111",
	"00111111",
	"00011110",
	"00000001",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"10000110",
	"11111011",
	"11111011",
	"11111011",
	"11111011",
	"11111111",
	"10000011",
	"11111011",
	"01111011",
	"10000110",
	"10000110",
	"10000110",
	"10001110",
	"01111010",
	"11111110",
	"10000110",
	"11111110",
	"11111110",
	"11111111",
	"11111100",
	"11110010",
	"10001110",
	"11111110",
	"11111111",
	"00000001",
	"00000001",
	"00000011",
	"00001111",
	"11111101",
	"11110001",
	"10000001",
	"01111110",
	"11111011",
	"11111011",
	"11111101",
	"11111101",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"10000110",
	"10000110",
	"10000011",
	"10000011",
	"10000001",
	"10000001",
	"11000001",
	"01111111",
	"00000000",
	"00000000",
	"11000000",
	"00110000",
	"00001000",
	"00000100",
	"00000010",
	"00000010",
	"00000000",
	"00000000",
	"11000000",
	"11110000",
	"11111000",
	"11111100",
	"11111110",
	"11111110",
	"00000000",
	"00000000",
	"00000011",
	"00001100",
	"00010000",
	"00100000",
	"01000000",
	"01000000",
	"00000000",
	"00000000",
	"00000011",
	"00001111",
	"00011111",
	"00111111",
	"01111111",
	"01111111",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00000010",
	"00000010",
	"00000010",
	"00000100",
	"00001100",
	"00111000",
	"11110000",
	"11100000",
	"11111110",
	"11111110",
	"11111110",
	"11111100",
	"11111100",
	"11111000",
	"11110000",
	"11100000",
	"01000000",
	"01000000",
	"01000000",
	"00100000",
	"00110000",
	"00011100",
	"00001111",
	"00001111",
	"01111111",
	"01111111",
	"01111111",
	"00111111",
	"00111111",
	"00011111",
	"00001111",
	"00001111",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00110000",
	"10100000",
	"01010000",
	"11110000",
	"11110000",
	"11110000",
	"11110000",
	"11110000",
	"11110000",
	"11100000",
	"11110000",
	"00001000",
	"00001010",
	"00001010",
	"00001010",
	"00001010",
	"00001100",
	"00000101",
	"00001010",
	"00001111",
	"00001111",
	"00001111",
	"00001111",
	"00001111",
	"00001111",
	"00000111",
	"00001111",
	"00000000",
	"10000010",
	"01000100",
	"01000100",
	"00111000",
	"00000000",
	"00000000",
	"00000000",
	"10000001",
	"10000011",
	"11000101",
	"11000101",
	"10111001",
	"10000001",
	"10000001",
	"10000001",
	"11000111",
	"00101000",
	"01111100",
	"01111100",
	"01111100",
	"01111100",
	"00101000",
	"11000111",
	"11000111",
	"11101111",
	"10000011",
	"10000011",
	"10000011",
	"10000011",
	"11101111",
	"11000111",
	"11111111",
	"11111111",
	"00011111",
	"00001111",
	"00001111",
	"00000111",
	"00000111",
	"00000111",
	"00000000",
	"00000000",
	"11100000",
	"11110000",
	"00110000",
	"11011000",
	"11011000",
	"11011000",
	"11111111",
	"11111111",
	"11111110",
	"11111100",
	"11111100",
	"11111001",
	"11111001",
	"11111001",
	"00000000",
	"00000000",
	"00000111",
	"00001111",
	"00001111",
	"00011111",
	"00011111",
	"00011111",
	"00000111",
	"00000111",
	"00000111",
	"00000111",
	"00000111",
	"11001111",
	"00001111",
	"00011111",
	"11011000",
	"11011000",
	"11011000",
	"11011000",
	"11011000",
	"11110000",
	"11110000",
	"11100000",
	"11111001",
	"11111001",
	"11111001",
	"11111001",
	"11111001",
	"11111100",
	"11111100",
	"11111110",
	"00011111",
	"00011111",
	"00011111",
	"00011111",
	"00011111",
	"00001111",
	"00001111",
	"00000111",
	"00000000",
	"00001110",
	"11111000",
	"00001000",
	"00001110",
	"11111110",
	"11111110",
	"11111110",
	"00000111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00000000",
	"11000000",
	"00011111",
	"00000000",
	"11000000",
	"11011111",
	"11011111",
	"11011111",
	"11100000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00111110",
	"11011110",
	"01101110",
	"10101110",
	"10101110",
	"11101110",
	"11101000",
	"11100110",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"01111111",
	"11111111",
	"11110111",
	"11011100",
	"11011111",
	"11011110",
	"11011111",
	"11011111",
	"11001111",
	"00011111",
	"11001111",
	"11111111",
	"11111011",
	"11110111",
	"11110101",
	"11110101",
	"11110110",
	"11110111",
	"11100111",
	"11110000",
	"11110000",
	"11111000",
	"11111000",
	"11111100",
	"00111100",
	"00011110",
	"01011110",
	"11111000",
	"11111000",
	"11111100",
	"11111100",
	"00001110",
	"11000110",
	"11100111",
	"10100111",
	"00011111",
	"00011111",
	"00111111",
	"00111111",
	"01111111",
	"01111100",
	"01111000",
	"11111010",
	"00001111",
	"00001111",
	"00011111",
	"00011111",
	"00110000",
	"00100011",
	"00100111",
	"01100101",
	"01101110",
	"01101110",
	"01101110",
	"00001110",
	"10111110",
	"00111110",
	"11111110",
	"11111110",
	"10010111",
	"10010111",
	"10010111",
	"11110111",
	"01000111",
	"11000111",
	"00001111",
	"11111111",
	"11110110",
	"11110110",
	"11110110",
	"11110000",
	"11111101",
	"11111100",
	"11111111",
	"11111111",
	"01101001",
	"01101001",
	"01101001",
	"01101111",
	"01100010",
	"01100011",
	"01110000",
	"01111111",
	"00111100",
	"01111110",
	"01111110",
	"11111111",
	"11111111",
	"11111111",
	"01000010",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01111110",
	"00111100",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00111100",
	"01000010",
	"10011001",
	"10000101",
	"10000101",
	"10011001",
	"01000010",
	"00111100",
	"00001111",
	"00000111",
	"00000111",
	"00000011",
	"00000011",
	"00000001",
	"00000001",
	"00000001",
	"11110000",
	"11111000",
	"11111000",
	"11111100",
	"11111100",
	"11111110",
	"11111110",
	"11111110",
	"11110000",
	"11100000",
	"11100000",
	"11000000",
	"11000000",
	"10000000",
	"10000000",
	"10000000",
	"00001111",
	"00011111",
	"00011111",
	"00111111",
	"00111111",
	"01111111",
	"01111111",
	"01111111",
	"00000001",
	"00000001",
	"00000011",
	"00000011",
	"00000111",
	"00011111",
	"01111111",
	"11111111",
	"11111110",
	"11111110",
	"11111100",
	"11111100",
	"11111100",
	"11111100",
	"11111000",
	"11111000",
	"11111111",
	"11111110",
	"11111000",
	"11100000",
	"11000000",
	"11000000",
	"10000000",
	"10000001",
	"01111111",
	"11111111",
	"11111111",
	"11111111",
	"00111111",
	"00111111",
	"01111111",
	"01111111",
	"00000001",
	"00000001",
	"00000001",
	"00000011",
	"00000011",
	"00000111",
	"00000111",
	"00001111",
	"11111110",
	"11111110",
	"11111110",
	"11111100",
	"11111100",
	"11111100",
	"11111100",
	"11111000",
	"10000000",
	"10000000",
	"10000000",
	"11000000",
	"11000000",
	"11100000",
	"11100000",
	"11110000",
	"01111111",
	"01111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"01111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111000",
	"11110000",
	"11110000",
	"11100000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"01111111",
	"00111111",
	"00111111",
	"00011111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"01111110",
	"01111110",
	"01111110",
	"01111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"10000000",
	"10000000",
	"10000000",
	"11000000",
	"11000000",
	"11100000",
	"11100000",
	"11110000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"01111111",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"01111111",
	"01111111",
	"01111111",
	"01111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111111",
	"11000000",
	"11000000",
	"11000000",
	"11000000",
	"11000000",
	"11000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00111111",
	"01111111",
	"01111111",
	"01111110",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"10000000",
	"10000000",
	"10000000",
	"11000000",
	"11100000",
	"11000000",
	"10000000",
	"10000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"01111111",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"01111110",
	"01111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111100",
	"11111100",
	"11111100",
	"11111100",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"01111110",
	"00111110",
	"00111110",
	"00011110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"01111111",
	"01111111",
	"11111111",
	"11111111",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"00000001",
	"00000001",
	"00000011",
	"00000011",
	"00000111",
	"00011111",
	"01111111",
	"11111111",
	"11111110",
	"11111110",
	"11111100",
	"11111100",
	"11111100",
	"11111100",
	"11111000",
	"11111000",
	"11111111",
	"11111110",
	"11111000",
	"11100000",
	"11000000",
	"11000000",
	"10000000",
	"10000001",
	"11111100",
	"11111101",
	"11111111",
	"11111111",
	"00111111",
	"00111111",
	"01111111",
	"01111111",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"11111110",
	"11111110",
	"01111110",
	"01111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"10000001",
	"01111110",
	"01111110",
	"01111110",
	"01111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"01111110",
	"00111100",
	"00111100",
	"00011000",
	"00011000",
	"00000000",
	"00000000",
	"00000000",
	"10000001",
	"11000011",
	"11000011",
	"11100111",
	"11100111",
	"11111111",
	"11111111",
	"11111111",
	"01001111",
	"01111111",
	"01111111",
	"11111111",
	"11111111",
	"11110111",
	"11101111",
	"00011111",
	"11110000",
	"11000010",
	"11011010",
	"11001010",
	"10001100",
	"10011000",
	"11110000",
	"11100000",
	"11111101",
	"01111101",
	"10111101",
	"11011110",
	"11011110",
	"11100000",
	"11001111",
	"10111111",
	"10000011",
	"11000011",
	"01100011",
	"00100001",
	"00111111",
	"00111111",
	"01110000",
	"01000000",
	"11111111",
	"11111111",
	"11111111",
	"11100110",
	"10011010",
	"01111001",
	"11111101",
	"11111101",
	"00001000",
	"00000100",
	"01000100",
	"01011101",
	"01100111",
	"10000111",
	"00000011",
	"00000011",
	"00000100",
	"01100111",
	"00101010",
	"01100100",
	"10000100",
	"01100000",
	"00101010",
	"01100100",
	"00000100",
	"01100101",
	"00101010",
	"01100100",
	"00000100",
	"01100011",
	"00101010",
	"01100100",
	"00000100",
	"01011001",
	"10000000",
	"10010010",
	"00000100",
	"10100101",
	"10010011",
	"01100010",
	"00000100",
	"10100001",
	"10000000",
	"00100010",
	"00000100",
	"01100001",
	"00101010",
	"00010010",
	"10001011",
	"00011011",
	"00011011",
	"01111011",
	"10001011",
	"00001011",
	"01011011",
	"01111011",
	"00000100",
	"01011101",
	"10010011",
	"01010010",
	"00000100",
	"01100101",
	"01010000",
	"00001011",
	"11011011",
	"10011011",
	"11011011",
	"00111011",
	"11011011",
	"11111011",
	"00000100",
	"01100111",
	"10001011",
	"00000100",
	"01100011",
	"01010000",
	"01001011",
	"11001011",
	"11011011",
	"11011011",
	"01011011",
	"11011011",
	"00000111",
	"10000100",
	"01100000",
	"01010000",
	"01101011",
	"11101011",
	"01010000",
	"00101011",
	"10101011",
	"00101011",
	"10011011",
	"11011011",
	"01000111",
	"00101011",
	"10000100",
	"01100100",
	"00101000",
	"00001011",
	"00010111",
	"10001011",
	"00001011",
	"10001011",
	"01101011",
	"11101011",
	"10000111",
	"01100100",
	"01101011",
	"10111011",
	"10000111",
	"10000111",
	"01111011",
	"10001011",
	"00001011",
	"10001011",
	"00001011",
	"10001011",
	"01100100",
	"10000100",
	"01111011",
	"10001011",
	"00011011",
	"00001011",
	"10001011",
	"01100100",
	"01111011",
	"10001011",
	"01000010",
	"11011011",
	"11011011",
	"01000010",
	"01100100",
	"11011011",
	"01000010",
	"11011011",
	"01100010",
	"00101000",
	"11011011",
	"01000010",
	"01000010",
	"11011011",
	"01000010",
	"11011011",
	"01100010",
	"11011011",
	"10000100",
	"00110110",
	"01110000",
	"11111011",
	"11011011",
	"11011011",
	"01000010",
	"11011011",
	"01000010",
	"11011011",
	"01000010",
	"01100100",
	"10000100",
	"01100110",
	"00100111",
	"10100111",
	"01100100",
	"10000100",
	"01100001",
	"00101000",
	"11011011",
	"11011011",
	"11011011",
	"01100100",
	"11011011",
	"11111011",
	"11011011",
	"11111011",
	"11011011",
	"11011011",
	"01100100",
	"11011011",
	"11000111",
	"11011011",
	"00000111",
	"11011011",
	"11011011",
	"01100111",
	"11011011",
	"01111011",
	"11000010",
	"11011011",
	"00000111",
	"11011011",
	"11011011",
	"11011011",
	"11011011",
	"01000010",
	"11011011",
	"11011011",
	"11011011",
	"00101011",
	"10011011",
	"01100100",
	"11000111",
	"01100100",
	"10000100",
	"01100101",
	"00101000",
	"11011011",
	"11011011",
	"11011011",
	"11100111",
	"10000100",
	"10100011",
	"01101000",
	"11111010",
	"10101001",
	"10101001",
	"10101001",
	"11011011",
	"10011011",
	"11011011",
	"11011011",
	"00101011",
	"10011011",
	"00101011",
	"10011011",
	"10101001",
	"01101001",
	"10101001",
	"10101001",
	"11101001",
	"00011001",
	"11101001",
	"00011001",
	"10101001",
	"10101001",
	"10101001",
	"10101001",
	"10101001",
	"11101001",
	"00011001",
	"00011110",
	"00010000",
	"10100000",
	"00100100",
	"11101000",
	"01001000",
	"11101000",
	"10111000",
	"01110000",
	"10101001",
	"01011110",
	"10000100",
	"10110111",
	"01110000",
	"11110011",
	"10000000",
	"10010000",
	"10011000",
	"10101000",
	"01010000",
	"01000100",
	"01110000",
	"11011000",
	"00100100",
	"00001000",
	"11101000",
	"10110000",
	"00011000",
	"01000100",
	"11010010",
	"10110000",
	"10000000",
	"00100100",
	"10011000",
	"10101000",
	"01010000",
	"01000100",
	"01110000",
	"11011000",
	"00100100",
	"00001000",
	"01010000",
	"01101000",
	"01110000",
	"01000100",
	"11010001",
	"10110000",
	"01000000",
	"00100100",
	"10011000",
	"00010100",
	"01000100",
	"01101111",
	"10000000",
	"00000000",
	"11000100",
	"10010011",
	"01010000",
	"01101000",
	"01110000",
	"01000100",
	"00110111",
	"00100000",
	"10111000",
	"00011000",
	"01010101",
	"11000100",
	"01010111",
	"00100000",
	"10011001",
	"01010101",
	"01010101",
	"01010101",
	"01101010",
	"10101010",
	"11000100",
	"01000111",
	"00100000",
	"10011001",
	"01010101",
	"01010101",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111000",
	"11111100",
	"11111100",
	"11111110",
	"11000000",
	"11110000",
	"11111000",
	"11111000",
	"00111000",
	"00100100",
	"01100100",
	"01100110",
	"00000000",
	"00000100",
	"00000110",
	"00000000",
	"00001111",
	"00111111",
	"01111111",
	"01111111",
	"00000111",
	"00000011",
	"00000001",
	"00111111",
	"00000001",
	"00000011",
	"00000000",
	"00000100",
	"11111110",
	"11111110",
	"11111000",
	"11100000",
	"00000000",
	"01111000",
	"11111100",
	"11111110",
	"00000110",
	"00001110",
	"00011000",
	"11100000",
	"11110000",
	"11111000",
	"11111100",
	"11111110",
	"00111111",
	"00111111",
	"00011111",
	"00000011",
	"01000011",
	"11100110",
	"11110100",
	"11101100",
	"00111111",
	"00111110",
	"00000000",
	"00000000",
	"00000111",
	"00001111",
	"00011111",
	"00011111",
	"11111110",
	"01111110",
	"00111111",
	"00001111",
	"00011111",
	"00011111",
	"00001111",
	"00001110",
	"11111110",
	"11111110",
	"11111111",
	"11111111",
	"11100000",
	"11100000",
	"11110000",
	"11110000",
	"11101100",
	"01101100",
	"00111010",
	"00000000",
	"00000000",
	"10000000",
	"11000000",
	"11111000",
	"10111111",
	"01111111",
	"00101101",
	"00011111",
	"00011111",
	"10011111",
	"11011111",
	"11111111",
	"00010000",
	"00100100",
	"11000111",
	"00001111",
	"00011111",
	"00001110",
	"00001110",
	"00011100",
	"11111000",
	"11111100",
	"11111111",
	"11111111",
	"00111111",
	"00001110",
	"00001110",
	"00011100",
	"11111000",
	"11111000",
	"11111000",
	"11111000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111111",
	"11111111",
	"11111111",
	"11111000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11110000",
	"11111000",
	"00000000",
	"00000000",
	"10000000",
	"11100000",
	"11110000",
	"11110000",
	"01110000",
	"01001000",
	"00000000",
	"00000000",
	"00000000",
	"00001000",
	"00001100",
	"00000000",
	"00011111",
	"01111111",
	"00000000",
	"00000000",
	"00001111",
	"00000111",
	"00000011",
	"01111111",
	"00000010",
	"00000110",
	"11111000",
	"11111100",
	"11111100",
	"11111000",
	"11100000",
	"00010000",
	"11101000",
	"11101000",
	"11001000",
	"11001100",
	"00001100",
	"00011000",
	"00100000",
	"11110000",
	"11111000",
	"11111000",
	"11111111",
	"11111111",
	"01111111",
	"01111111",
	"00111111",
	"00000111",
	"00000010",
	"00000101",
	"00000000",
	"00001000",
	"01111110",
	"01111100",
	"00000000",
	"00000000",
	"00000011",
	"00000111",
	"11101100",
	"11100100",
	"11000100",
	"11000000",
	"10000000",
	"00000000",
	"00000000",
	"00000000",
	"11111100",
	"11111100",
	"11111100",
	"11111000",
	"11111000",
	"11111000",
	"11111000",
	"11111000",
	"00110011",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00001110",
	"00000000",
	"00010000",
	"00001111",
	"00001111",
	"00001111",
	"00011111",
	"00011111",
	"00011111",
	"00011111",
	"00011111",
	"00001111",
	"00001111",
	"00001111",
	"00001111",
	"00001111",
	"00000011",
	"00000001",
	"00000000",
	"11111111",
	"11111111",
	"11111111",
	"01111111",
	"00001111",
	"00000011",
	"00000001",
	"00000000",
	"00001000",
	"00000110",
	"00000001",
	"00000000",
	"00011110",
	"00011110",
	"01111110",
	"01111110",
	"00111111",
	"00111111",
	"00011111",
	"00011110",
	"00011110",
	"00011110",
	"01111110",
	"01111110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111000",
	"11111100",
	"11111100",
	"00000000",
	"11000000",
	"11110000",
	"11111000",
	"11111000",
	"00111000",
	"00100100",
	"01100100",
	"00000000",
	"00000000",
	"00000100",
	"00000110",
	"00000000",
	"00001111",
	"00111111",
	"01111111",
	"00000000",
	"00000111",
	"00000011",
	"00000001",
	"00111111",
	"00000001",
	"00000011",
	"00000000",
	"11111110",
	"11111110",
	"11111100",
	"11111000",
	"00000000",
	"01101000",
	"11110100",
	"11110100",
	"01100110",
	"00000110",
	"00001100",
	"00011000",
	"11110000",
	"11111000",
	"11111100",
	"11111100",
	"01111111",
	"00111111",
	"00111111",
	"00011111",
	"00000011",
	"00000110",
	"00000100",
	"00001100",
	"00000100",
	"00111111",
	"00111110",
	"00000000",
	"00000000",
	"00000111",
	"00000111",
	"00001111",
	"11110100",
	"11110100",
	"11110100",
	"11110000",
	"11100000",
	"11000000",
	"00000000",
	"00000000",
	"11111100",
	"11111100",
	"11111100",
	"11111100",
	"11111100",
	"11111100",
	"11111100",
	"11111000",
	"00001000",
	"00001111",
	"00001111",
	"00001111",
	"00001111",
	"00000111",
	"00000011",
	"00000111",
	"00001111",
	"00001001",
	"00000000",
	"00010000",
	"00110000",
	"00111000",
	"00111111",
	"00011111",
	"10000000",
	"11000000",
	"10000000",
	"00100000",
	"11100000",
	"11110000",
	"11110000",
	"11000000",
	"11110000",
	"11110000",
	"11100000",
	"11100000",
	"11100000",
	"11110000",
	"11110000",
	"11000000",
	"00011111",
	"00001111",
	"00000111",
	"00001110",
	"00001101",
	"00000001",
	"00000111",
	"00000111",
	"00011111",
	"00001111",
	"00000111",
	"00001111",
	"00001101",
	"00000001",
	"00000111",
	"00000111",
	"00000000",
	"00001100",
	"00001110",
	"11111110",
	"11111111",
	"11111111",
	"11101111",
	"11001111",
	"11000000",
	"11111100",
	"11111110",
	"10011000",
	"10010000",
	"10010000",
	"00010100",
	"00111010",
	"00000000",
	"00011000",
	"00001000",
	"00000000",
	"00011111",
	"00011111",
	"01111111",
	"11111111",
	"00011111",
	"00000111",
	"00000111",
	"00111111",
	"01100100",
	"00001100",
	"00000001",
	"00001000",
	"11100111",
	"11110000",
	"11110000",
	"11111000",
	"11111000",
	"11111000",
	"11110000",
	"11100000",
	"01111100",
	"01111000",
	"11111100",
	"00011100",
	"00001100",
	"00001100",
	"00000000",
	"01011100",
	"11111111",
	"01111111",
	"00111111",
	"01100011",
	"01110001",
	"01110111",
	"11111111",
	"11111111",
	"00011110",
	"01111000",
	"00000001",
	"01111111",
	"01111110",
	"01111110",
	"11111110",
	"11111110",
	"11000000",
	"00000000",
	"00000000",
	"01110000",
	"11100000",
	"11111100",
	"11111100",
	"11111100",
	"00111100",
	"11111100",
	"11111000",
	"11110000",
	"11100000",
	"11111100",
	"10000100",
	"00000100",
	"11111111",
	"11111110",
	"11111100",
	"01110000",
	"00000011",
	"00000011",
	"00000111",
	"00000111",
	"11111111",
	"11111111",
	"11111111",
	"01111111",
	"01111111",
	"01111111",
	"00111111",
	"00001110",
	"00000000",
	"00000001",
	"00010011",
	"01111111",
	"11111110",
	"11111100",
	"01111000",
	"01110000",
	"11110000",
	"11111001",
	"11110011",
	"11111111",
	"11111110",
	"11111100",
	"01111000",
	"01110000",
	"00000111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000100",
	"00000011",
	"00000001",
	"00000001",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111000",
	"11111100",
	"00000000",
	"00000000",
	"11000000",
	"11110000",
	"11111000",
	"11111000",
	"00111000",
	"00100100",
	"01110000",
	"11111000",
	"11111000",
	"11111000",
	"11111000",
	"11000000",
	"11111111",
	"11111111",
	"00000000",
	"00100000",
	"01100111",
	"00000111",
	"11111111",
	"11111111",
	"11110001",
	"11000001",
	"11111100",
	"11111100",
	"11111110",
	"11111110",
	"11111000",
	"00000000",
	"01111110",
	"11111111",
	"01100100",
	"01100100",
	"00000110",
	"00011110",
	"00011000",
	"11110000",
	"11111110",
	"11111111",
	"11111111",
	"11111111",
	"01111111",
	"01111111",
	"01111111",
	"01111011",
	"00111010",
	"00110110",
	"10000000",
	"10000100",
	"01111111",
	"01011110",
	"01100000",
	"01111111",
	"00111111",
	"00111111",
	"11111111",
	"11111111",
	"01111111",
	"00111111",
	"00011111",
	"00001101",
	"00000110",
	"00000000",
	"11111111",
	"11110011",
	"11100001",
	"11100000",
	"11100000",
	"11110000",
	"11111000",
	"11111000",
	"00010100",
	"00001100",
	"00011000",
	"00000010",
	"00000000",
	"10000000",
	"11000000",
	"11110000",
	"00011111",
	"00011111",
	"00001111",
	"00011101",
	"00011111",
	"10011111",
	"11011111",
	"11111111",
	"00001000",
	"00110111",
	"11000111",
	"00000111",
	"00000111",
	"00000111",
	"00000011",
	"00000001",
	"11111000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"01111111",
	"00000011",
	"00000001",
	"11110000",
	"11110000",
	"11110000",
	"11110000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111111",
	"11111111",
	"11111111",
	"11111100",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111000",
	"11111100",
	"11111100",
	"11111000",
	"11100000",
	"10010000",
	"11001000",
	"11101000",
	"11001000",
	"11001100",
	"00001100",
	"00011000",
	"00100000",
	"11110000",
	"11111000",
	"11111000",
	"11111111",
	"11111111",
	"01111111",
	"11111111",
	"01111111",
	"00111111",
	"00011111",
	"00000111",
	"00000000",
	"00001000",
	"01111110",
	"00001100",
	"00000111",
	"00001111",
	"00001111",
	"00000111",
	"11101000",
	"11101000",
	"11000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111000",
	"11111000",
	"11110000",
	"11110000",
	"11110000",
	"11111000",
	"11111000",
	"11111000",
	"00001011",
	"00001001",
	"00011000",
	"00010000",
	"00000010",
	"00000000",
	"00000000",
	"00000000",
	"00001111",
	"00001111",
	"00011111",
	"00011111",
	"00011101",
	"00011111",
	"00011111",
	"00011111",
	"00001100",
	"00001111",
	"00001111",
	"10001111",
	"01101111",
	"01100011",
	"00100001",
	"00000000",
	"11111100",
	"11111111",
	"11111111",
	"11111111",
	"01101111",
	"01100011",
	"00100001",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00001111",
	"00000111",
	"00000001",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111000",
	"11111000",
	"11111100",
	"01111100",
	"00111110",
	"00011110",
	"00001111",
	"00000111",
	"11111000",
	"11111000",
	"11111100",
	"11111100",
	"11111000",
	"11110000",
	"11110000",
	"11111000",
	"00001101",
	"00001001",
	"00011000",
	"00010000",
	"00000010",
	"00000000",
	"00000000",
	"00000000",
	"00001111",
	"00001111",
	"00011111",
	"00011111",
	"00011101",
	"00011111",
	"00011111",
	"00001111",
	"00000011",
	"00000111",
	"00111111",
	"01111111",
	"11111111",
	"11111110",
	"11000000",
	"00000000",
	"00000111",
	"00001111",
	"00001111",
	"00001111",
	"00001111",
	"00001111",
	"00011111",
	"00001111",
	"00000000",
	"00000000",
	"00001000",
	"00011100",
	"01111100",
	"00111100",
	"00011100",
	"00011000",
	"11111000",
	"11111000",
	"11111000",
	"11111100",
	"01111100",
	"00111100",
	"00011100",
	"00011000",
	"00000000",
	"00000000",
	"00000000",
	"11100000",
	"11110000",
	"11110000",
	"11110000",
	"11000000",
	"00000000",
	"11000000",
	"11100000",
	"11100000",
	"01010000",
	"11010000",
	"00110000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00001111",
	"00111111",
	"01111111",
	"00111111",
	"00011111",
	"00000000",
	"00000111",
	"00111111",
	"00000100",
	"00000100",
	"00001000",
	"00111100",
	"00000000",
	"11100000",
	"11110000",
	"11011000",
	"00011000",
	"00001000",
	"00001100",
	"10000100",
	"10000000",
	"11100000",
	"11100000",
	"11100000",
	"11111000",
	"11111000",
	"01111100",
	"10000100",
	"10000000",
	"00010101",
	"00111111",
	"00011111",
	"00000000",
	"00000000",
	"00000000",
	"00000011",
	"00000111",
	"00000111",
	"00000111",
	"00000111",
	"00001111",
	"00001111",
	"00000111",
	"00000011",
	"00000111",
	"00000000",
	"00000000",
	"11110000",
	"11111000",
	"11111000",
	"11111000",
	"11100000",
	"00111100",
	"11100000",
	"11110000",
	"01110000",
	"00101000",
	"01101000",
	"00011000",
	"00000000",
	"11111100",
	"00000000",
	"00000000",
	"00000111",
	"00011111",
	"00111111",
	"00011111",
	"00001111",
	"00000011",
	"00000011",
	"00011111",
	"00000010",
	"00000010",
	"00000100",
	"00011110",
	"00000000",
	"00000011",
	"00111111",
	"10110111",
	"00000011",
	"00000000",
	"00000000",
	"00000110",
	"00001110",
	"00011100",
	"11111100",
	"01110000",
	"11110000",
	"11111000",
	"11111100",
	"00111110",
	"00001110",
	"00011100",
	"01111110",
	"01111000",
	"00100000",
	"00110000",
	"00110000",
	"00110000",
	"00000000",
	"00000000",
	"00001111",
	"00011111",
	"00100111",
	"00111111",
	"00111111",
	"00111110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11110000",
	"11111000",
	"11111000",
	"11111000",
	"11100000",
	"10110000",
	"11100000",
	"11110000",
	"01110000",
	"00101000",
	"01101000",
	"00011000",
	"00000000",
	"11110000",
	"01111000",
	"00111000",
	"01111000",
	"11110000",
	"11100000",
	"00000000",
	"11100000",
	"11100000",
	"11111000",
	"11111000",
	"11111000",
	"00111000",
	"00110000",
	"11100000",
	"11100000",
	"11100000",
	"00000110",
	"00001001",
	"00000000",
	"00000001",
	"00000000",
	"00000111",
	"00001111",
	"00000001",
	"00000111",
	"00000110",
	"00001111",
	"00001110",
	"00000111",
	"00000111",
	"00001111",
	"00000001",
	"00000000",
	"00001000",
	"11111100",
	"11111110",
	"11111110",
	"11111100",
	"11000000",
	"11110000",
	"11100000",
	"11111000",
	"11111100",
	"01001000",
	"11001000",
	"00010000",
	"11111000",
	"10001100",
	"00000000",
	"00000000",
	"00000111",
	"00011111",
	"00111111",
	"00011111",
	"00001101",
	"00011100",
	"00000011",
	"00001111",
	"00000010",
	"00000000",
	"00001100",
	"00011000",
	"00000011",
	"00011111",
	"11111000",
	"11100000",
	"00000000",
	"01110000",
	"11110000",
	"11001010",
	"00111110",
	"00111100",
	"10001100",
	"10011100",
	"11111000",
	"11111000",
	"11110000",
	"11111010",
	"01111110",
	"00111100",
	"00011111",
	"00011111",
	"00001111",
	"00000000",
	"00000000",
	"00000001",
	"00000000",
	"00000000",
	"00011111",
	"00011111",
	"00001111",
	"00000111",
	"00000111",
	"00000011",
	"00000000",
	"00000000",
	"11100000",
	"11100000",
	"11000000",
	"11101111",
	"11111111",
	"11111111",
	"01111111",
	"00111111",
	"00000000",
	"00000111",
	"00111111",
	"11100100",
	"11100100",
	"10001000",
	"01111100",
	"00100000",
	"01111100",
	"11111110",
	"11111111",
	"01000111",
	"00001010",
	"00011100",
	"00001110",
	"00000010",
	"11111100",
	"11111110",
	"11111100",
	"11110000",
	"11111000",
	"11111100",
	"11111110",
	"11110010",
	"00010111",
	"10001110",
	"10000000",
	"11010010",
	"11000000",
	"11000000",
	"00000000",
	"00000000",
	"00011111",
	"10011111",
	"10011111",
	"11101101",
	"11111111",
	"11111111",
	"00000111",
	"00000000",
	"10100000",
	"11000000",
	"10000000",
	"00001100",
	"00001100",
	"00001100",
	"01100100",
	"00100000",
	"11100000",
	"11100000",
	"11110000",
	"11111100",
	"11111100",
	"11111100",
	"01100100",
	"00100000",
	"01111111",
	"00111111",
	"00000111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00001111",
	"00001111",
	"00001111",
	"00000111",
	"00000011",
	"00000000",
	"00000000",
	"00000000",
	"10100000",
	"11000000",
	"10000000",
	"00001000",
	"00001100",
	"00110000",
	"00111000",
	"00011000",
	"11100000",
	"11100000",
	"11110000",
	"11111000",
	"11111100",
	"11110000",
	"00111000",
	"00011000",
	"00000011",
	"00000111",
	"00001111",
	"00011110",
	"00011000",
	"00010000",
	"00000000",
	"00000000",
	"00000111",
	"00000111",
	"00000111",
	"00000111",
	"00000011",
	"00000001",
	"00000000",
	"00000000",
	"11100000",
	"11110000",
	"01111100",
	"00111110",
	"00001100",
	"00110000",
	"00111000",
	"00011000",
	"11100000",
	"11110000",
	"11111000",
	"11110000",
	"11111100",
	"11110000",
	"00111000",
	"00011000",
	"00000110",
	"00000110",
	"00000110",
	"00000001",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000111",
	"00000111",
	"00000111",
	"00000010",
	"00000011",
	"00000001",
	"00000000",
	"00000000",
	"11001110",
	"11001111",
	"00001111",
	"00101111",
	"00001111",
	"00001111",
	"00001110",
	"00000110",
	"11111110",
	"11111111",
	"11111111",
	"11011111",
	"11110000",
	"11110000",
	"11110000",
	"11111000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00111100",
	"00111100",
	"00111111",
	"00111111",
	"11111100",
	"01111110",
	"00111110",
	"00111110",
	"00111100",
	"00111100",
	"00111111",
	"00111111",
	"11111110",
	"11111110",
	"11111000",
	"11100000",
	"11010000",
	"11011000",
	"11011100",
	"11011110",
	"00000110",
	"00001110",
	"00011000",
	"00010000",
	"11110000",
	"11111000",
	"11111100",
	"11111110",
	"00111111",
	"00111111",
	"00011111",
	"00000111",
	"00001011",
	"00011011",
	"00111011",
	"01111011",
	"00111111",
	"00111110",
	"00000000",
	"00000100",
	"00001111",
	"00011111",
	"00111111",
	"01111111",
	"00100011",
	"00000111",
	"00000111",
	"00000010",
	"00000000",
	"00111100",
	"00111100",
	"00111110",
	"11010000",
	"11110000",
	"11111000",
	"01111000",
	"00111100",
	"00111100",
	"00111100",
	"00111110",
	"10111000",
	"00111100",
	"01011100",
	"00011100",
	"00001100",
	"00000000",
	"00111000",
	"00111100",
	"11111000",
	"11111100",
	"10110000",
	"11100000",
	"11110000",
	"01110000",
	"00111000",
	"00111100",
	"01000100",
	"10101010",
	"10101010",
	"10101010",
	"10101010",
	"10101010",
	"11101110",
	"01000100",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11100000",
	"11111000",
	"11111111",
	"11100000",
	"11111000",
	"11110000",
	"01100000",
	"00000000",
	"00000000",
	"11110011",
	"11100000",
	"11111110",
	"00000000",
	"00000000",
	"00000000",
	"11111100",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11011111",
	"01101110",
	"00000000",
	"00000000",
	"00111100",
	"00111111",
	"01111111",
	"00000111",
	"00000000",
	"00000000",
	"00000100",
	"00011111",
	"11111111",
	"11000011",
	"10111111",
	"01111111",
	"00001111",
	"00000010",
	"00000010",
	"00000111",
	"00000010",
	"11111100",
	"01111100",
	"01111100",
	"00001100",
	"00011100",
	"00000010",
	"00000111",
	"00000010",
	"00000010",
	"10000010",
	"10000010",
	"11110010",
	"11100010",
	"00000000",
	"00000000",
	"00000000",
	"00011111",
	"00011111",
	"00011111",
	"00011000",
	"00011100",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000111",
	"00000011",
	"00111100",
	"10011100",
	"11011100",
	"11111100",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11000010",
	"01100010",
	"00100010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00011110",
	"00011100",
	"00011101",
	"00011111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000001",
	"00000011",
	"00000010",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111100",
	"11111100",
	"11110000",
	"11101110",
	"11101110",
	"11101111",
	"11101111",
	"11101111",
	"10001100",
	"00001100",
	"00011100",
	"00111110",
	"11111110",
	"11111111",
	"11111111",
	"11011111",
	"11111111",
	"01111111",
	"01111111",
	"01111111",
	"01011111",
	"01011111",
	"11001111",
	"11100111",
	"00001000",
	"01111110",
	"01111100",
	"00000000",
	"01111000",
	"01111111",
	"11111111",
	"11111111",
	"00001111",
	"00011111",
	"00111111",
	"00111110",
	"00011110",
	"00011100",
	"00111100",
	"00111111",
	"11111111",
	"11111111",
	"11000111",
	"11000011",
	"11100001",
	"00010010",
	"00111100",
	"00111111",
	"11111111",
	"00000000",
	"11000011",
	"10000001",
	"10000001",
	"11000011",
	"11111111",
	"00000000",
	"00000000",
	"11111111",
	"11000011",
	"11000001",
	"11000001",
	"11111111",
	"11111111",
	"11111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111000",
	"11111000",
	"11110000",
	"11100000",
	"10000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11010000",
	"11111000",
	"11111000",
	"01111000",
	"01111100",
	"00110000",
	"00100000",
	"00001111",
	"11011111",
	"11111111",
	"11111111",
	"01111111",
	"01111100",
	"00110000",
	"00100000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111000",
	"11111000",
	"11110000",
	"11110000",
	"11100000",
	"00000000",
	"00000000",
	"00000000",
	"11000000",
	"11110000",
	"11110000",
	"11110000",
	"11110000",
	"00000000",
	"00000000",
	"00000000",
	"11011111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00011000",
	"00111100",
	"01111110",
	"01101110",
	"11011111",
	"11011111",
	"11011111",
	"00000000",
	"00011000",
	"00111100",
	"01111110",
	"01110110",
	"11111011",
	"11111011",
	"11111011",
	"00000000",
	"00001000",
	"00001000",
	"00000100",
	"00000100",
	"00000100",
	"00000100",
	"00000100",
	"00000000",
	"00011000",
	"00011000",
	"00111100",
	"00111100",
	"00111100",
	"00111100",
	"00111000",
	"00000000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00000000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00000000",
	"00000000",
	"00001000",
	"00001000",
	"00011100",
	"00011100",
	"00011100",
	"00011100",
	"00011100",
	"00000000",
	"00010000",
	"00010000",
	"00100000",
	"00100000",
	"00100000",
	"00100000",
	"00100000",
	"00000000",
	"00011000",
	"00111100",
	"01110000",
	"01110000",
	"00100000",
	"00000000",
	"00000000",
	"00111100",
	"01111110",
	"11101110",
	"11011111",
	"11111001",
	"11111010",
	"01110001",
	"00000100",
	"00000000",
	"00000000",
	"00100000",
	"01100000",
	"01111000",
	"00111100",
	"00011000",
	"00000000",
	"00111010",
	"01110100",
	"11110001",
	"11111100",
	"11011110",
	"11101110",
	"01111110",
	"00111100",
	"00000000",
	"00000000",
	"10000000",
	"01010000",
	"11101000",
	"11110000",
	"11110100",
	"11111000",
	"11001000",
	"11110010",
	"11111100",
	"11111101",
	"11111100",
	"01011110",
	"00011111",
	"00011111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"10100000",
	"11100000",
	"11110000",
	"11100000",
	"00000000",
	"00010000",
	"10100000",
	"11110000",
	"11110100",
	"10111000",
	"00111000",
	"00111100",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"10000000",
	"11000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01000000",
	"11010000",
	"11100000",
	"11110000",
	"00000000",
	"00000110",
	"00001111",
	"00011111",
	"00111110",
	"01111100",
	"01111110",
	"11111110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00010000",
	"00100000",
	"00100000",
	"11111100",
	"11111010",
	"11111110",
	"01111100",
	"01110000",
	"01010000",
	"10001010",
	"00000100",
	"01000000",
	"01000000",
	"01000000",
	"10100000",
	"10001110",
	"11111110",
	"11111110",
	"11111110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01110000",
	"11111000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00100000",
	"11111100",
	"11111110",
	"11111110",
	"01111111",
	"00110111",
	"01010011",
	"10001010",
	"00000100",
	"01000000",
	"01000000",
	"00000000",
	"10000000",
	"11001000",
	"11111100",
	"11111110",
	"11111110",
	"00000000",
	"00000010",
	"11000110",
	"11101110",
	"00111110",
	"00011100",
	"00011111",
	"00100111",
	"00000000",
	"00000010",
	"00000110",
	"00001110",
	"11001110",
	"11100100",
	"11110000",
	"11111000",
	"00000000",
	"00000000",
	"11000000",
	"11100000",
	"00110000",
	"00011000",
	"00011111",
	"00100111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11000000",
	"11100000",
	"11110000",
	"11111000",
	"11000000",
	"00100010",
	"00010100",
	"00001000",
	"00010000",
	"00100000",
	"11000000",
	"00100000",
	"11111110",
	"11111110",
	"11111100",
	"11111100",
	"11111000",
	"11111000",
	"11110000",
	"11100000",
	"11000000",
	"11100000",
	"11110000",
	"11111000",
	"11100100",
	"11011110",
	"00011110",
	"11011111",
	"11000000",
	"11100000",
	"11110000",
	"11111000",
	"11111100",
	"11101110",
	"11101110",
	"10101111",
	"00000011",
	"00000111",
	"00001111",
	"00011111",
	"00100111",
	"01111011",
	"01111000",
	"11111011",
	"00000011",
	"00000111",
	"00001111",
	"00011111",
	"00111111",
	"01110111",
	"01110111",
	"11110101",
	"11111111",
	"11111111",
	"11111110",
	"11110000",
	"11110000",
	"11100000",
	"11000000",
	"00000000",
	"10001111",
	"11111111",
	"00011110",
	"00000000",
	"00000000",
	"00011000",
	"00111000",
	"01110000",
	"11111111",
	"11111111",
	"01111111",
	"00001111",
	"00001111",
	"00000011",
	"00000001",
	"00000000",
	"11110001",
	"11111111",
	"01111000",
	"00000000",
	"00110000",
	"01111100",
	"01111110",
	"00111110",
	"00000000",
	"00000000",
	"00011000",
	"00100100",
	"00100100",
	"00011000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00111100",
	"01111110",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"01111110",
	"00111100",
	"00000000",
	"01000000",
	"10000010",
	"10000010",
	"10000110",
	"11001100",
	"01100000",
	"00111100",
	"11000000",
	"11100000",
	"11110000",
	"11111000",
	"11111100",
	"11000110",
	"10000010",
	"10000011",
	"11000000",
	"11100000",
	"11110000",
	"11111000",
	"11111100",
	"11111110",
	"11111110",
	"11111111",
	"00000011",
	"00000001",
	"00000000",
	"00000000",
	"00110001",
	"01111111",
	"01111111",
	"11001111",
	"00000011",
	"00000111",
	"00001111",
	"00011111",
	"00111111",
	"01111111",
	"01111111",
	"11111111",
	"10000011",
	"11000111",
	"11111111",
	"11100010",
	"11110000",
	"11110000",
	"11110000",
	"11100000",
	"11111111",
	"11111111",
	"11111111",
	"00011110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"10001111",
	"10011111",
	"11111111",
	"01000111",
	"00001111",
	"00001111",
	"00001111",
	"00000111",
	"11111111",
	"11111111",
	"11111111",
	"01111000",
	"00000000",
	"00000100",
	"00000100",
	"00000010",
	"01101000",
	"11111000",
	"00000000",
	"00000000",
	"10100000",
	"10110000",
	"11111100",
	"11111000",
	"01101000",
	"11111000",
	"11111100",
	"11111110",
	"10111100",
	"10111000",
	"11111100",
	"11111000",
	"00000001",
	"00000001",
	"00000000",
	"00000000",
	"00000000",
	"00000101",
	"00000101",
	"00000111",
	"00000001",
	"00000001",
	"00000011",
	"00000111",
	"00001111",
	"00001111",
	"00001111",
	"00011111",
	"00000000",
	"00100000",
	"01110010",
	"00110001",
	"00110000",
	"11111110",
	"11111111",
	"11111111",
	"00111100",
	"01011111",
	"10001101",
	"01001110",
	"01001111",
	"11011011",
	"11111011",
	"11111010",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"10000000",
	"10000000",
	"00000000",
	"00000000",
	"00000000",
	"10000000",
	"10000000",
	"10000000",
	"01100000",
	"01111000",
	"11111111",
	"11111110",
	"11111100",
	"11111000",
	"11110000",
	"11100000",
	"11000000",
	"10000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111111",
	"11000001",
	"10010100",
	"10110110",
	"10100010",
	"10001000",
	"10000000",
	"11100011",
	"00000000",
	"00111110",
	"01101011",
	"01001001",
	"01011101",
	"01110111",
	"01111111",
	"00011100",
	"00010000",
	"00010000",
	"01000000",
	"11111000",
	"01000100",
	"01000000",
	"01000000",
	"00000000",
	"00000000",
	"10101000",
	"11111100",
	"01000110",
	"11111010",
	"11111111",
	"11111001",
	"10111110",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00010000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00001000",
	"01111000",
	"00001000",
	"00001010",
	"00001000",
	"00010000",
	"00000000",
	"00000000",
	"11110100",
	"01111000",
	"11110100",
	"11110100",
	"11110100",
	"10101000",
	"10110000",
	"01110000",
	"00000000",
	"00000000",
	"00000000",
	"01111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00111000",
	"01010100",
	"11101110",
	"01110111",
	"10111011",
	"01010101",
	"00101110",
	"00010100",
	"00111000",
	"01111100",
	"11111110",
	"11111111",
	"11111111",
	"01111111",
	"00111110",
	"00011100",
	"11111111",
	"01111111",
	"01111111",
	"00000000",
	"11110111",
	"11110111",
	"11110111",
	"00000000",
	"00000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"01111111",
	"01111111",
	"01111111",
	"00000000",
	"11110111",
	"11110111",
	"11110111",
	"00000000",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00000000",
	"11111110",
	"11111010",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"11111111",
	"00011101",
	"01111001",
	"00000001",
	"00000011",
	"00000111",
	"00001111",
	"00011111",
	"00111110",
	"00010110",
	"01110010",
	"00000111",
	"00000111",
	"00000111",
	"00001111",
	"00011111",
	"00111111",
	"00000000",
	"11000100",
	"11101010",
	"11110010",
	"11101010",
	"11100100",
	"11000011",
	"10000100",
	"11111100",
	"00111010",
	"10011100",
	"11011100",
	"11011101",
	"10011111",
	"00111111",
	"01111111",
	"00000000",
	"00001100",
	"00001110",
	"00001110",
	"00001111",
	"00000111",
	"00000011",
	"00000000",
	"00000011",
	"00001111",
	"00001111",
	"00001111",
	"00001111",
	"00000111",
	"00000011",
	"00000000",
	"11001000",
	"11110000",
	"01111000",
	"00001111",
	"00111111",
	"00011111",
	"00001111",
	"00000111",
	"01111111",
	"00111111",
	"10000110",
	"11110000",
	"11111111",
	"01111111",
	"00001111",
	"00000111",
	"01111101",
	"00001001",
	"00000001",
	"00000011",
	"00000011",
	"00000001",
	"00000000",
	"00000000",
	"01110110",
	"00000010",
	"00000111",
	"00000111",
	"00000111",
	"00000111",
	"00000111",
	"00000011",
	"10000000",
	"10000000",
	"11000000",
	"11000000",
	"11100000",
	"11111110",
	"10111110",
	"10111100",
	"10000000",
	"10000000",
	"11000000",
	"11000000",
	"11100000",
	"11111110",
	"11111110",
	"11111100",
	"01100000",
	"00100000",
	"00001100",
	"11000100",
	"01100000",
	"00100110",
	"00000110",
	"00000000",
	"01100000",
	"11100000",
	"11111100",
	"00111100",
	"10011000",
	"11011110",
	"11111110",
	"11111100",
	"00000000",
	"00000110",
	"00000110",
	"00000000",
	"00000100",
	"00001100",
	"00100000",
	"01100000",
	"11111100",
	"11111110",
	"11111110",
	"11111000",
	"11111100",
	"11111100",
	"11100000",
	"01100000",
	"00000000",
	"10000000",
	"10000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11000000",
	"11100000",
	"11110000",
	"11110000",
	"11110000",
	"11110000",
	"11100000",
	"11000000",
	"01111111",
	"11111111",
	"11111111",
	"00000010",
	"10000000",
	"11000000",
	"11000000",
	"11000000",
	"00011111",
	"00011111",
	"00011111",
	"00000101",
	"10000111",
	"11111111",
	"11111111",
	"11111111",
	"10000000",
	"10000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11110000",
	"11110000",
	"11110000",
	"11111000",
	"11111000",
	"11111000",
	"11110000",
	"11100000",
	"00000111",
	"01111111",
	"11111111",
	"11111110",
	"11000000",
	"01000000",
	"00000000",
	"00000000",
	"00000111",
	"00011111",
	"00011111",
	"00011111",
	"11111111",
	"01111111",
	"00001111",
	"00000011",
	"10000000",
	"10110000",
	"00010000",
	"00000000",
	"01101100",
	"00110100",
	"00010000",
	"00000110",
	"10000000",
	"11110000",
	"11110000",
	"11111000",
	"10011100",
	"11001100",
	"11101100",
	"11111110",
	"00000110",
	"00000000",
	"00000100",
	"00001100",
	"00000000",
	"00010000",
	"10110000",
	"10000000",
	"11111110",
	"11111100",
	"11111100",
	"11111100",
	"11111000",
	"11110000",
	"11110000",
	"10000000",
	"10000000",
	"10000000",
	"11000000",
	"11000010",
	"11100110",
	"11101110",
	"11011110",
	"00011110",
	"00000000",
	"00000000",
	"11000000",
	"11000000",
	"11100010",
	"11100110",
	"11101110",
	"11101110",
	"00000000",
	"00000000",
	"00000001",
	"00100001",
	"00110011",
	"00111011",
	"00111101",
	"00111100",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00010001",
	"00011001",
	"00011111",
	"00001111",
	"11001100",
	"11100000",
	"11100000",
	"11000111",
	"00011100",
	"11111100",
	"00111000",
	"00110000",
	"01111110",
	"11111110",
	"11111111",
	"11111000",
	"11100000",
	"00001100",
	"00111000",
	"00110000",
	"00011001",
	"11100011",
	"00010011",
	"01001001",
	"00001100",
	"00011111",
	"00001110",
	"00000110",
	"01111110",
	"00011100",
	"01101111",
	"10110111",
	"11111011",
	"00011100",
	"00001110",
	"00000110",
	"00000000",
	"10000000",
	"10000000",
	"11000000",
	"11000010",
	"11100110",
	"11101110",
	"11011110",
	"00000000",
	"00000000",
	"00000000",
	"11000000",
	"11000000",
	"11100010",
	"11100110",
	"11101110",
	"00000000",
	"00000000",
	"00000000",
	"00000001",
	"00100001",
	"00110011",
	"00111011",
	"00111101",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00010001",
	"00011001",
	"00011111",
	"00011110",
	"11001100",
	"11100000",
	"11100000",
	"11000111",
	"00011100",
	"11111110",
	"00001111",
	"11101110",
	"01111110",
	"11111110",
	"11111111",
	"11111000",
	"11100000",
	"00001110",
	"00001111",
	"00111100",
	"00011001",
	"11100011",
	"00010011",
	"01001001",
	"00001100",
	"00011111",
	"00111100",
	"00001111",
	"01111110",
	"00011100",
	"01101111",
	"10110111",
	"11111011",
	"00011100",
	"00111100",
	"00000000",
	"00001000",
	"11111110",
	"11111110",
	"11111110",
	"11111000",
	"11110000",
	"11110000",
	"11000000",
	"11100000",
	"01010000",
	"01011000",
	"00111000",
	"01111000",
	"11010000",
	"00010000",
	"11000000",
	"11001100",
	"10011100",
	"01011100",
	"00011100",
	"00011000",
	"00000000",
	"00000000",
	"00111000",
	"11111100",
	"11111100",
	"10111100",
	"11111100",
	"11111000",
	"00000000",
	"00000000",
	"00001000",
	"00011100",
	"00111100",
	"00101110",
	"01101110",
	"01101110",
	"01111110",
	"10111110",
	"00000000",
	"00000000",
	"00100000",
	"00110010",
	"01110010",
	"01110010",
	"01100010",
	"11110110",
	"00000000",
	"00000000",
	"10001000",
	"01010000",
	"00101100",
	"01010100",
	"10001010",
	"00000100",
	"00000000",
	"11111000",
	"11111100",
	"11111100",
	"11110010",
	"11111010",
	"11111110",
	"11111110",
	"11111110",
	"11100110",
	"11000110",
	"00001110",
	"00011100",
	"01111100",
	"00111110",
	"00011101",
	"11111110",
	"11100110",
	"11000101",
	"00001101",
	"00011011",
	"01111011",
	"00111011",
	"00010011",
	"10001010",
	"01010000",
	"00100000",
	"01010111",
	"10011110",
	"11111110",
	"00001110",
	"10011100",
	"11111110",
	"11111110",
	"11111110",
	"11111000",
	"11100010",
	"00001110",
	"00001110",
	"10011100",
	"00011010",
	"00011100",
	"00001000",
	"00001100",
	"00001111",
	"00001111",
	"00000111",
	"00000011",
	"00010111",
	"00010111",
	"00000111",
	"00000011",
	"00001000",
	"00001110",
	"00000111",
	"00000011",
	"00000000",
	"00010000",
	"00111000",
	"00111100",
	"01011110",
	"01011110",
	"01011110",
	"01111110",
	"00000000",
	"00000000",
	"00000000",
	"00000100",
	"01100110",
	"01100110",
	"01100110",
	"01000110",
	"00000000",
	"00000000",
	"00000000",
	"10001000",
	"01010000",
	"00101100",
	"01010100",
	"10001010",
	"00000000",
	"00000000",
	"11111000",
	"11111100",
	"11111110",
	"11110010",
	"11111010",
	"11111110",
	"11111110",
	"10111110",
	"11111100",
	"11101100",
	"11001100",
	"11011100",
	"01011100",
	"00011110",
	"11101110",
	"11111110",
	"11111100",
	"11101101",
	"11001101",
	"11011011",
	"01011011",
	"00011011",
	"00000100",
	"10001010",
	"01010000",
	"00100000",
	"01010111",
	"10011100",
	"11111110",
	"00001111",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111000",
	"11100000",
	"00001110",
	"00001111",
	"00111101",
	"00011010",
	"00011100",
	"00001000",
	"00001100",
	"00011111",
	"00111111",
	"01111100",
	"00110011",
	"00010111",
	"00010111",
	"00000111",
	"00000011",
	"00011000",
	"00111110",
	"01111100",
	"00000000",
	"00000000",
	"00000000",
	"01100000",
	"01110000",
	"00110000",
	"00000000",
	"00000000",
	"11000000",
	"11110000",
	"11111000",
	"11111100",
	"11011100",
	"11111100",
	"11111110",
	"11111110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11110000",
	"00011000",
	"00000001",
	"00001111",
	"00011111",
	"00111111",
	"01111111",
	"01111111",
	"11111111",
	"01111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00011111",
	"01111100",
	"11011100",
	"00011000",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111111",
	"11110000",
	"11000000",
	"00000000",
	"00001000",
	"00101000",
	"00001000",
	"00001000",
	"00011100",
	"00011110",
	"00011111",
	"00001100",
	"01111111",
	"11011111",
	"11111111",
	"11111111",
	"01101111",
	"00000111",
	"00000011",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01100000",
	"01110000",
	"00110000",
	"00000000",
	"00000000",
	"11000000",
	"11110000",
	"11111000",
	"11111100",
	"11011100",
	"11111100",
	"11111110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11110000",
	"00000000",
	"00000011",
	"00001111",
	"00011111",
	"00111111",
	"01111111",
	"01111111",
	"11111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00011111",
	"01111110",
	"11001111",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111111",
	"11110000",
	"11000000",
	"00011000",
	"00001000",
	"00101000",
	"00001000",
	"00001000",
	"00011100",
	"00111110",
	"01111011",
	"01111111",
	"01111111",
	"11011111",
	"11111111",
	"11111111",
	"01101111",
	"00000111",
	"00000011",
	"00000000",
	"10110000",
	"01111000",
	"01111000",
	"01111000",
	"11111000",
	"11110000",
	"11100000",
	"00000000",
	"10000000",
	"10000000",
	"10000000",
	"10000000",
	"00000000",
	"00000000",
	"00010000",
	"00011110",
	"00001111",
	"00000000",
	"01011000",
	"11111100",
	"10101100",
	"10101100",
	"11111100",
	"00011110",
	"00001111",
	"00011111",
	"00100111",
	"00000011",
	"01010011",
	"01010011",
	"00000011",
	"00000000",
	"00000000",
	"00000001",
	"00000111",
	"00000111",
	"00001110",
	"11001110",
	"10000100",
	"11110000",
	"11111000",
	"11111001",
	"11111111",
	"11111111",
	"11111110",
	"00101110",
	"00000100",
	"01011000",
	"11100000",
	"00110000",
	"00011000",
	"00011110",
	"01111111",
	"00111111",
	"00001111",
	"00100111",
	"11111111",
	"01111111",
	"00111111",
	"00111001",
	"01111000",
	"00000000",
	"00000000",
	"00000000",
	"10000000",
	"01000000",
	"00000000",
	"00011100",
	"00111110",
	"01111110",
	"11111100",
	"00000000",
	"10000000",
	"11000000",
	"11000000",
	"11100000",
	"11000000",
	"10000000",
	"00000000",
	"11111100",
	"00000010",
	"00000110",
	"00000110",
	"00000100",
	"00001100",
	"11001000",
	"10000000",
	"00000000",
	"11111010",
	"11111110",
	"11111110",
	"11111100",
	"11111100",
	"00101000",
	"00000000",
	"00000011",
	"00000111",
	"00001100",
	"00001011",
	"00001011",
	"00001011",
	"00001011",
	"00000000",
	"00000011",
	"00000111",
	"00001111",
	"00001100",
	"00011100",
	"00111100",
	"00111100",
	"00111111",
	"11100000",
	"11110000",
	"01000000",
	"10111000",
	"11111000",
	"01011000",
	"01011000",
	"01000000",
	"11100000",
	"11110000",
	"11111000",
	"01000100",
	"00000100",
	"10100100",
	"10100100",
	"11111000",
	"00011100",
	"00111110",
	"00111111",
	"00111111",
	"00111111",
	"01111111",
	"01111101",
	"01111101",
	"01111111",
	"01111111",
	"01111110",
	"01011100",
	"01000000",
	"10000000",
	"10000010",
	"10000010",
	"00111000",
	"01111100",
	"11111100",
	"11111100",
	"11111100",
	"11111110",
	"10111110",
	"10111110",
	"11111000",
	"11111100",
	"01111110",
	"00111010",
	"00000010",
	"00000001",
	"01000001",
	"01000001",
	"10111110",
	"11111110",
	"11111010",
	"11011100",
	"00111100",
	"11111100",
	"01111000",
	"00000000",
	"01000001",
	"00000001",
	"00000101",
	"00100010",
	"11000010",
	"00000010",
	"10000100",
	"01111000",
	"00111000",
	"01111100",
	"11111100",
	"11111000",
	"11111100",
	"11111110",
	"10111110",
	"10111110",
	"00111000",
	"11111100",
	"01111100",
	"00111100",
	"00000010",
	"00000001",
	"01000001",
	"01000001",
	"00000000",
	"00000000",
	"00000000",
	"00000110",
	"01000110",
	"10100110",
	"11111100",
	"11111000",
	"00000000",
	"00000000",
	"00000001",
	"00000001",
	"01001001",
	"10111001",
	"11100011",
	"11110111",
	"00001110",
	"00111100",
	"00111100",
	"00011000",
	"00000000",
	"00000000",
	"01000000",
	"11100000",
	"00000000",
	"11000100",
	"11001100",
	"11111100",
	"11111100",
	"11111110",
	"11111110",
	"11111110",
	"11110011",
	"01011110",
	"01011010",
	"00001000",
	"00000000",
	"00000000",
	"00000011",
	"00000001",
	"01111111",
	"00011111",
	"00000101",
	"00000000",
	"00000000",
	"00000000",
	"00000001",
	"00000001",
	"10100001",
	"00100001",
	"01100001",
	"01100011",
	"11100111",
	"11001110",
	"11001110",
	"10000111",
	"01111110",
	"11111110",
	"10111110",
	"11111100",
	"01111000",
	"11110001",
	"11110001",
	"10011000",
	"00000001",
	"01110010",
	"11101110",
	"11001111",
	"11011111",
	"10011111",
	"01011111",
	"00011110",
	"00000111",
	"01110000",
	"11001110",
	"11001111",
	"10011111",
	"10011111",
	"00011111",
	"00001110",
	"10001000",
	"10011100",
	"10111110",
	"10011100",
	"00000000",
	"00000000",
	"00000111",
	"11100111",
	"01110000",
	"01100110",
	"01000111",
	"01101111",
	"11111111",
	"11111111",
	"11111000",
	"00011001",
	"00000000",
	"00000000",
	"11100000",
	"11100000",
	"01101000",
	"00001000",
	"00000000",
	"00011100",
	"00000000",
	"00000000",
	"00000000",
	"00100000",
	"11110000",
	"11110000",
	"11111000",
	"11100000",
	"11110011",
	"11111000",
	"11101000",
	"00001000",
	"11001100",
	"00001100",
	"00001100",
	"00000100",
	"11001111",
	"11100111",
	"01110111",
	"00110111",
	"10110011",
	"11110011",
	"11110011",
	"11111011",
	"00011100",
	"00001100",
	"00000010",
	"11100011",
	"11100000",
	"01100110",
	"00000111",
	"00110110",
	"11100100",
	"11111100",
	"11111100",
	"00011110",
	"00111100",
	"11111000",
	"11111000",
	"11001110",
	"00000110",
	"00000011",
	"00000001",
	"00100000",
	"01111001",
	"11111111",
	"00001111",
	"00011111",
	"11111001",
	"01111100",
	"00111110",
	"00111111",
	"00011111",
	"00011111",
	"00000011",
	"00000010",
	"00100100",
	"10000000",
	"11100000",
	"01111111",
	"11111111",
	"11111110",
	"11111100",
	"11111110",
	"11111110",
	"01111110",
	"00011110",
	"10000000",
	"11100000",
	"11111000",
	"00111100",
	"00111110",
	"11110011",
	"01011110",
	"01010000",
	"01111111",
	"00111111",
	"00000000",
	"00000000",
	"00000000",
	"00111111",
	"00011111",
	"00000101",
	"01111111",
	"00111111",
	"00001111",
	"00000001",
	"00000000",
	"10100001",
	"01100001",
	"11000001",
	"11000011",
	"10000111",
	"00001110",
	"00001110",
	"00000111",
	"01111110",
	"11111110",
	"11111110",
	"11111100",
	"11111000",
	"11110001",
	"11110001",
	"00011000",
	"00000110",
	"00000011",
	"00000001",
	"00000000",
	"00011001",
	"00111111",
	"01111111",
	"11111111",
	"11111001",
	"01111100",
	"00111110",
	"00011111",
	"00011111",
	"00111100",
	"00011000",
	"00011111",
	"00100100",
	"00000000",
	"11100000",
	"01111111",
	"11111111",
	"11111110",
	"11111111",
	"11000000",
	"11111110",
	"11111110",
	"00011110",
	"10000000",
	"11100000",
	"11001000",
	"10001111",
	"11000000",
	"11000000",
	"11110000",
	"11000100",
	"01000110",
	"00100110",
	"00111100",
	"00111000",
	"01111000",
	"00000000",
	"00000000",
	"00111000",
	"10111000",
	"11011000",
	"11000011",
	"11000111",
	"10000111",
	"11111000",
	"10111100",
	"10110110",
	"11110010",
	"01110111",
	"11001111",
	"00000100",
	"11000000",
	"00000111",
	"10110011",
	"10111000",
	"11110010",
	"01110111",
	"11111111",
	"11111100",
	"11111100",
	"11100000",
	"11100000",
	"11111000",
	"11111100",
	"11110000",
	"11100010",
	"11000000",
	"00000000",
	"11111100",
	"11111100",
	"00000000",
	"00000000",
	"00001110",
	"00011101",
	"00111111",
	"00111111",
	"00000000",
	"00000000",
	"11000000",
	"11100000",
	"11110000",
	"11110000",
	"11111000",
	"11111000",
	"11100000",
	"11110000",
	"11111000",
	"11111100",
	"01111100",
	"00111110",
	"00011110",
	"00011110",
	"00000000",
	"11000100",
	"11101010",
	"11110010",
	"11101010",
	"11110100",
	"11111011",
	"10000100",
	"11111100",
	"00111010",
	"10011100",
	"11011100",
	"11111101",
	"11111111",
	"01111111",
	"01111111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000001",
	"00000001",
	"00000000",
	"00000000",
	"00000011",
	"00000011",
	"00000001",
	"00000001",
	"00000001",
	"00000001",
	"00000000",
	"00000000",
	"11000100",
	"11110000",
	"01111000",
	"00001111",
	"00111000",
	"11111100",
	"11111000",
	"01111000",
	"01111111",
	"00111111",
	"10000110",
	"11110000",
	"11111110",
	"11111100",
	"11111000",
	"01111000",
	"00000000",
	"00000001",
	"00011000",
	"00001100",
	"00101100",
	"01111111",
	"01111111",
	"01111111",
	"00001111",
	"00011110",
	"00100111",
	"00010011",
	"00110011",
	"01111101",
	"01111101",
	"01111100",
	"00000000",
	"00000000",
	"10000000",
	"00100000",
	"01100000",
	"01100000",
	"11100000",
	"11100000",
	"00000000",
	"10000000",
	"00000000",
	"11100000",
	"11100000",
	"11100000",
	"11100000",
	"11111000",
	"11110000",
	"11111100",
	"11111110",
	"00011111",
	"00011111",
	"11111110",
	"11111100",
	"11110000",
	"00000000",
	"00000000",
	"11110000",
	"11111100",
	"11111100",
	"11110000",
	"00000000",
	"00000000",
	"11111000",
	"11111000",
	"11111000",
	"11010000",
	"10000000",
	"10000000",
	"00000000",
	"00000000",
	"00011110",
	"00111110",
	"01111110",
	"11111110",
	"11111100",
	"11111100",
	"11011000",
	"10010000",
	"11000000",
	"11111000",
	"11111100",
	"11111100",
	"00011110",
	"00000000",
	"11000000",
	"11111111",
	"00110000",
	"00000000",
	"00000000",
	"00000000",
	"11100000",
	"11111110",
	"00111110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"10000000",
	"10000111",
	"10001110",
	"10011110",
	"10111100",
	"10111100",
	"11111000",
	"11000000",
	"11000100",
	"11100100",
	"11111000",
	"11100000",
	"11110000",
	"11111000",
	"11111110",
	"11111100",
	"11111100",
	"11111100",
	"11111000",
	"11011000",
	"01101100",
	"00001100",
	"11111110",
	"11111100",
	"00000111",
	"00000001",
	"00000001",
	"00000010",
	"00000111",
	"00000111",
	"00000111",
	"00000011",
	"00011111",
	"00011111",
	"00011111",
	"00011101",
	"00011000",
	"00011011",
	"00011011",
	"00011101",
	"11000000",
	"11100000",
	"11110000",
	"11111000",
	"11111100",
	"11111110",
	"11111111",
	"11111000",
	"10000000",
	"01000000",
	"00100000",
	"00100000",
	"00010000",
	"00010000",
	"00001000",
	"00001000",
	"11111000",
	"00001000",
	"00110000",
	"01001000",
	"01001000",
	"00110100",
	"11111100",
	"11111100",
	"00000000",
	"11110000",
	"11001000",
	"10110000",
	"10110000",
	"11001000",
	"00110000",
	"00000100",
	"11101100",
	"01101100",
	"01101100",
	"01101100",
	"01101000",
	"01101000",
	"01001000",
	"01000000",
	"00000000",
	"00100100",
	"00000000",
	"00100100",
	"00000000",
	"00100000",
	"00000000",
	"00000000",
	"00001000",
	"01111110",
	"11111111",
	"11111111",
	"01101111",
	"01101110",
	"01011100",
	"01011000",
	"11110000",
	"10000010",
	"00000000",
	"00010001",
	"00000000",
	"00100010",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00011100",
	"00100000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00011100",
	"00111110",
	"01111111",
	"01111111",
	"11011100",
	"11000000",
	"11000000",
	"11000000",
	"00000000",
	"00000000",
	"00000000",
	"00011100",
	"00000010",
	"00000000",
	"00000000",
	"00000000",
	"11000000",
	"11001100",
	"11011110",
	"11111110",
	"11111111",
	"11011111",
	"11000000",
	"11000000",
	"00111111",
	"00000101",
	"00000001",
	"00000001",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00111011",
	"00000011",
	"00000111",
	"00000111",
	"00000111",
	"00000111",
	"00000111",
	"00000011",
	"11100000",
	"11100100",
	"11101010",
	"11110010",
	"11101010",
	"11100100",
	"10000011",
	"10000100",
	"11111100",
	"11111010",
	"11111100",
	"11111100",
	"11011101",
	"00011111",
	"01111111",
	"01111111",
	"10111000",
	"11110000",
	"11110000",
	"11111000",
	"11111000",
	"01111000",
	"00011100",
	"00001100",
	"11111000",
	"11110000",
	"11110000",
	"11111000",
	"11111000",
	"01111000",
	"00011100",
	"00001100",
	"00000000",
	"00000000",
	"00011100",
	"00001000",
	"00110010",
	"00011000",
	"01100001",
	"00100100",
	"00000000",
	"00000100",
	"00000110",
	"00000110",
	"00001110",
	"00001111",
	"00011111",
	"00011111",
	"00000000",
	"01000010",
	"01010000",
	"00000010",
	"00001000",
	"01000000",
	"00010000",
	"01000000",
	"00011111",
	"00111111",
	"00111111",
	"01111110",
	"01111110",
	"01111100",
	"11111000",
	"11100000",
	"00000000",
	"00000000",
	"00000001",
	"00000010",
	"00010000",
	"00110000",
	"01010000",
	"00100001",
	"00000000",
	"00000011",
	"00001110",
	"00011101",
	"00101111",
	"01001111",
	"10101111",
	"11011110",
	"00000000",
	"00000000",
	"11110011",
	"00000100",
	"00000100",
	"00000100",
	"01100100",
	"01110100",
	"00000000",
	"11111011",
	"00001000",
	"11111111",
	"11111011",
	"11111111",
	"11111111",
	"10011111",
	"00000111",
	"00000111",
	"00000011",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11111000",
	"11111000",
	"01111100",
	"00111111",
	"00011111",
	"00001111",
	"00000011",
	"00000000",
	"11110100",
	"11000100",
	"10000100",
	"00000100",
	"00000100",
	"00000000",
	"00000000",
	"00000000",
	"00011111",
	"00111111",
	"01111111",
	"11111111",
	"11111111",
	"11111011",
	"11111011",
	"00000000",
	"10000011",
	"10001101",
	"10011010",
	"10110110",
	"10101100",
	"11011100",
	"11111000",
	"11000000",
	"10000011",
	"10001111",
	"10011110",
	"10111110",
	"10111100",
	"11111100",
	"11111000",
	"11000000",
	"00000000",
	"01000000",
	"00000000",
	"00010000",
	"01000000",
	"00000000",
	"00010100",
	"00000000",
	"01000000",
	"01100000",
	"01110000",
	"01110000",
	"01111000",
	"01111000",
	"01111100",
	"01111100",
	"00100000",
	"00001000",
	"01000000",
	"00001000",
	"00100000",
	"00000000",
	"01010000",
	"00000000",
	"01111100",
	"01111100",
	"01111100",
	"01111100",
	"01111000",
	"01111000",
	"01110000",
	"01000000",
	"10000011",
	"10001101",
	"10011010",
	"10110110",
	"10101100",
	"11011100",
	"11111000",
	"11000000",
	"10000011",
	"10001111",
	"10011110",
	"10111110",
	"10111100",
	"11111100",
	"11111000",
	"11000000",
	"00000000",
	"11110000",
	"11111000",
	"11111111",
	"00111111",
	"11000110",
	"11111000",
	"11000000",
	"00111110",
	"00000000",
	"00000000",
	"11111111",
	"11000011",
	"11111110",
	"11111000",
	"11000000",
	"00000000",
	"00000000",
	"01111111",
	"01100011",
	"01100011",
	"01111111",
	"00000000",
	"00000000",
	"11111111",
	"11111111",
	"00111110",
	"00000000",
	"00000000",
	"00111110",
	"11111111",
	"11111111",
	"00000000",
	"00000000",
	"01100000",
	"01100000",
	"00110000",
	"00011000",
	"00001110",
	"00000110",
	"11111111",
	"11111111",
	"00000000",
	"00100000",
	"00110000",
	"00011000",
	"00001100",
	"00000000",
	"00000000",
	"00000000",
	"01100000",
	"01100000",
	"00100000",
	"00100000",
	"00010000",
	"00010000",
	"11111111",
	"11111111",
	"00000000",
	"00100000",
	"00100000",
	"00100000",
	"00010000",
	"00010000",
	"00010000",
	"00001000",
	"00001100",
	"00001100",
	"00001100",
	"00001100",
	"00001000",
	"00010000",
	"00010000",
	"00001000",
	"00001000",
	"00000000",
	"00000000",
	"00001000",
	"00001000",
	"00010000",
	"00000000",
	"00000000",
	"10000000",
	"11000000",
	"10000000",
	"00000000",
	"00000000",
	"00000000",
	"11111110",
	"11111100",
	"11111100",
	"01111100",
	"11111000",
	"11110000",
	"11000000",
	"00000000",
	"11000000",
	"01110000",
	"00011111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"11000000",
	"11110000",
	"11111111",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"11111110",
	"01000100",
	"10100110",
	"10100100",
	"10100100",
	"10100100",
	"10100100",
	"11101110",
	"01001110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01000110",
	"10101001",
	"10101000",
	"10100100",
	"10100010",
	"10100001",
	"11101111",
	"01001111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01000101",
	"10100101",
	"10100101",
	"10100101",
	"10101111",
	"10101111",
	"11100100",
	"01000100",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01001111",
	"10100001",
	"10100001",
	"10100111",
	"10101000",
	"10101000",
	"11101111",
	"01000111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01000110",
	"10101001",
	"10101010",
	"10100110",
	"10101101",
	"10101001",
	"11101001",
	"01000110",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000100",
	"00001010",
	"00001010",
	"00001010",
	"00001010",
	"00001010",
	"00001110",
	"00000100",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01100110",
	"01100111",
	"01100110",
	"01100110",
	"01100110",
	"11100110",
	"11001111",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"01111010",
	"10011010",
	"10011010",
	"10011010",
	"01111010",
	"00011011",
	"00011001",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00100000",
	"00010000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00111110",
	"00011100",
	"00000000"
);

begin

dir_int_img <= to_integer(unsigned(dir_tabla_patrones));

P_img: process (clk)
begin
	if clk'event and clk='1' then
		dato_tabla_patrones <= title(dir_int_img);
	end if;
end process;

end behavioral;	
